//출처 : https://verilogguide.readthedocs.io/en/latest/verilog/designs.html#read-only-memory-rom

module ROM(
    input wire clk,
	input wire En,
    input wire  [13:0] addr,
    output reg signed [25:0] data1,
	output reg signed [25:0] data2,
	output reg signed [25:0] data3,
	output reg signed [25:0] data4
);

//ROM[0]?�� ?���?? : 16bit(?�� ?��그널?�� ?���??) * 4(4개의 ?��그널) 
// 각각?�� ?��그널?�� �?? 1000sample?�� ?��?���??�?? addr??  16비트�?? ?��?��(0~39999 < 0~65536) 

reg signed [25:0] ROM1[0:127];
reg signed [25:0] ROM2[0:127];
reg signed [25:0] ROM3[0:127];
reg signed [25:0] ROM4[0:127];
reg [6:0] cnt;

always @(posedge clk) begin
	if(!En) begin
		cnt<=0;
        data1<=0;
        data2<=0;
        data3<=0;
        data4<=0;

ROM1[0]<=-26'd12648; ROM2[0]<=-26'd10090; ROM3[0]<=-26'd46841; ROM4[0]<=-26'd29163;
ROM1[1]<=-26'd33679; ROM2[1]<=-26'd28067; ROM3[1]<=-26'd108968; ROM4[1]<=-26'd81697;
ROM1[2]<=-26'd30550; ROM2[2]<=-26'd24343; ROM3[2]<=-26'd93964; ROM4[2]<=-26'd80254;
ROM1[3]<=-26'd38879; ROM2[3]<=-26'd37267; ROM3[3]<=-26'd116594; ROM4[3]<=-26'd83223;
ROM1[4]<=-26'd43361; ROM2[4]<=-26'd43540; ROM3[4]<=-26'd119035; ROM4[4]<=-26'd91934;
ROM1[5]<=-26'd37302; ROM2[5]<=-26'd35397; ROM3[5]<=-26'd108666; ROM4[5]<=-26'd82744;
ROM1[6]<=-26'd35384; ROM2[6]<=-26'd30262; ROM3[6]<=-26'd98720; ROM4[6]<=-26'd91519;
ROM1[7]<=-26'd35061; ROM2[7]<=-26'd31834; ROM3[7]<=-26'd100315; ROM4[7]<=-26'd83473;
ROM1[8]<=-26'd42381; ROM2[8]<=-26'd41718; ROM3[8]<=-26'd111240; ROM4[8]<=-26'd95343;
ROM1[9]<=-26'd33003; ROM2[9]<=-26'd32672; ROM3[9]<=-26'd98195; ROM4[9]<=-26'd67998;
ROM1[10]<=-26'd41836; ROM2[10]<=-26'd38827; ROM3[10]<=-26'd101211; ROM4[10]<=-26'd106131;
ROM1[11]<=-26'd12294; ROM2[11]<=-26'd4004; ROM3[11]<=-26'd58622; ROM4[11]<=-26'd41210;
ROM1[12]<=26'd9241; ROM2[12]<=26'd19505; ROM3[12]<=-26'd30174; ROM4[12]<=26'd13514;
ROM1[13]<=-26'd32851; ROM2[13]<=-26'd28921; ROM3[13]<=-26'd88842; ROM4[13]<=-26'd83892;
ROM1[14]<=-26'd31868; ROM2[14]<=-26'd28628; ROM3[14]<=-26'd87250; ROM4[14]<=-26'd78992;
ROM1[15]<=-26'd40860; ROM2[15]<=-26'd38267; ROM3[15]<=-26'd94691; ROM4[15]<=-26'd104624;
ROM1[16]<=-26'd33562; ROM2[16]<=-26'd33114; ROM3[16]<=-26'd87196; ROM4[16]<=-26'd75831;
ROM1[17]<=-26'd29953; ROM2[17]<=-26'd28945; ROM3[17]<=-26'd81721; ROM4[17]<=-26'd67720;
ROM1[18]<=-26'd30483; ROM2[18]<=-26'd29355; ROM3[18]<=-26'd82808; ROM4[18]<=-26'd69386;
ROM1[19]<=-26'd39491; ROM2[19]<=-26'd39967; ROM3[19]<=-26'd95801; ROM4[19]<=-26'd89152;
ROM1[20]<=-26'd35325; ROM2[20]<=-26'd34299; ROM3[20]<=-26'd84215; ROM4[20]<=-26'd85193;
ROM1[21]<=-26'd42093; ROM2[21]<=-26'd46213; ROM3[21]<=-26'd98560; ROM4[21]<=-26'd84921;
ROM1[22]<=-26'd34938; ROM2[22]<=-26'd39892; ROM3[22]<=-26'd92605; ROM4[22]<=-26'd60086;
ROM1[23]<=-26'd38936; ROM2[23]<=-26'd47465; ROM3[23]<=-26'd102774; ROM4[23]<=-26'd57306;
ROM1[24]<=-26'd42370; ROM2[24]<=-26'd49184; ROM3[24]<=-26'd104917; ROM4[24]<=-26'd73755;
ROM1[25]<=-26'd38512; ROM2[25]<=-26'd46447; ROM3[25]<=-26'd100226; ROM4[25]<=-26'd58886;
ROM1[26]<=-26'd45508; ROM2[26]<=-26'd58856; ROM3[26]<=-26'd117438; ROM4[26]<=-26'd57106;
ROM1[27]<=-26'd44684; ROM2[27]<=-26'd56143; ROM3[27]<=-26'd112808; ROM4[27]<=-26'd62603;
ROM1[28]<=-26'd39524; ROM2[28]<=-26'd49974; ROM3[28]<=-26'd104617; ROM4[28]<=-26'd51850;
ROM1[29]<=-26'd55628; ROM2[29]<=-26'd77337; ROM3[29]<=-26'd139485; ROM4[29]<=-26'd54124;
ROM1[30]<=-26'd59097; ROM2[30]<=-26'd81866; ROM3[30]<=-26'd143697; ROM4[30]<=-26'd60662;
ROM1[31]<=-26'd49799; ROM2[31]<=-26'd68354; ROM3[31]<=-26'd124440; ROM4[31]<=-26'd51384;
ROM1[32]<=-26'd52368; ROM2[32]<=-26'd71144; ROM3[32]<=-26'd125510; ROM4[32]<=-26'd59076;
ROM1[33]<=-26'd32179; ROM2[33]<=-26'd44593; ROM3[33]<=-26'd90770; ROM4[33]<=-26'd26421;
ROM1[34]<=-26'd62341; ROM2[34]<=-26'd84912; ROM3[34]<=-26'd145489; ROM4[34]<=-26'd71581;
ROM1[35]<=-26'd59114; ROM2[35]<=-26'd81536; ROM3[35]<=-26'd146808; ROM4[35]<=-26'd60091;
ROM1[36]<=-26'd75758; ROM2[36]<=-26'd96387; ROM3[36]<=-26'd157050; ROM4[36]<=-26'd119035;
ROM1[37]<=26'd15029; ROM2[37]<=26'd8816; ROM3[37]<=-26'd28172; ROM4[37]<=26'd87442;
ROM1[38]<=26'd69611; ROM2[38]<=26'd68830; ROM3[38]<=26'd43309; ROM4[38]<=26'd225083;
ROM1[39]<=-26'd39450; ROM2[39]<=-26'd50561; ROM3[39]<=-26'd93356; ROM4[39]<=-26'd54737;
ROM1[40]<=-26'd25517; ROM2[40]<=-26'd30806; ROM3[40]<=-26'd66923; ROM4[40]<=-26'd38133;
ROM1[41]<=-26'd49151; ROM2[41]<=-26'd65324; ROM3[41]<=-26'd111553; ROM4[41]<=-26'd63190;
ROM1[42]<=-26'd39418; ROM2[42]<=-26'd55756; ROM3[42]<=-26'd99534; ROM4[42]<=-26'd34625;
ROM1[43]<=-26'd36971; ROM2[43]<=-26'd51015; ROM3[43]<=-26'd86631; ROM4[43]<=-26'd40016;
ROM1[44]<=-26'd25349; ROM2[44]<=-26'd34930; ROM3[44]<=-26'd63865; ROM4[44]<=-26'd25275;
ROM1[45]<=-26'd37231; ROM2[45]<=-26'd51285; ROM3[45]<=-26'd86399; ROM4[45]<=-26'd41114;
ROM1[46]<=-26'd33762; ROM2[46]<=-26'd45324; ROM3[46]<=-26'd78957; ROM4[46]<=-26'd40852;
ROM1[47]<=-26'd35272; ROM2[47]<=-26'd50387; ROM3[47]<=-26'd85545; ROM4[47]<=-26'd31358;
ROM1[48]<=-26'd32426; ROM2[48]<=-26'd49404; ROM3[48]<=-26'd84084; ROM4[48]<=-26'd16138;
ROM1[49]<=-26'd33260; ROM2[49]<=-26'd49447; ROM3[49]<=-26'd86246; ROM4[49]<=-26'd20617;
ROM1[50]<=-26'd25270; ROM2[50]<=-26'd35955; ROM3[50]<=-26'd63746; ROM4[50]<=-26'd21853;
ROM1[51]<=-26'd27788; ROM2[51]<=-26'd38662; ROM3[51]<=-26'd66187; ROM4[51]<=-26'd28901;
ROM1[52]<=-26'd30248; ROM2[52]<=-26'd42106; ROM3[52]<=-26'd72570; ROM4[52]<=-26'd31193;
ROM1[53]<=-26'd28933; ROM2[53]<=-26'd39235; ROM3[53]<=-26'd66276; ROM4[53]<=-26'd34862;
ROM1[54]<=-26'd25416; ROM2[54]<=-26'd35455; ROM3[54]<=-26'd57659; ROM4[54]<=-26'd27774;
ROM1[55]<=-26'd17138; ROM2[55]<=-26'd22594; ROM3[55]<=-26'd34324; ROM4[55]<=-26'd25423;
ROM1[56]<=-26'd20733; ROM2[56]<=-26'd30262; ROM3[56]<=-26'd47719; ROM4[56]<=-26'd18128;
ROM1[57]<=-26'd22911; ROM2[57]<=-26'd35420; ROM3[57]<=-26'd56096; ROM4[57]<=-26'd11922;
ROM1[58]<=-26'd20375; ROM2[58]<=-26'd32136; ROM3[58]<=-26'd50513; ROM4[58]<=-26'd8314;
ROM1[59]<=-26'd25203; ROM2[59]<=-26'd41243; ROM3[59]<=-26'd65990; ROM4[59]<=-26'd3597;
ROM1[60]<=-26'd13159; ROM2[60]<=-26'd21992; ROM3[60]<=-26'd38620; ROM4[60]<=26'd1429;
ROM1[61]<=-26'd9737; ROM2[61]<=-26'd16107; ROM3[61]<=-26'd27261; ROM4[61]<=-26'd297;
ROM1[62]<=-26'd13102; ROM2[62]<=-26'd17474; ROM3[62]<=-26'd31156; ROM4[62]<=-26'd16626;
ROM1[63]<=-26'd11613; ROM2[63]<=-26'd16170; ROM3[63]<=-26'd27122; ROM4[63]<=-26'd12831;
ROM1[64]<=-26'd7151; ROM2[64]<=-26'd11308; ROM3[64]<=-26'd17001; ROM4[64]<=-26'd3566;
ROM1[65]<=-26'd13066; ROM2[65]<=-26'd17866; ROM3[65]<=-26'd25483; ROM4[65]<=-26'd17922;
ROM1[66]<=-26'd2682; ROM2[66]<=-26'd2821; ROM3[66]<=-26'd2734; ROM4[66]<=-26'd8068;
ROM1[67]<=-26'd2974; ROM2[67]<=-26'd2171; ROM3[67]<=26'd413; ROM4[67]<=-26'd13692;
ROM1[68]<=26'd3069; ROM2[68]<=26'd2630; ROM3[68]<=26'd6065; ROM4[68]<=26'd8715;
ROM1[69]<=26'd7616; ROM2[69]<=26'd9505; ROM3[69]<=26'd15534; ROM4[69]<=26'd12378;
ROM1[70]<=26'd2738; ROM2[70]<=26'd2662; ROM3[70]<=26'd7147; ROM4[70]<=26'd5937;
ROM1[71]<=26'd12285; ROM2[71]<=26'd14117; ROM3[71]<=26'd25655; ROM4[71]<=26'd23958;
ROM1[72]<=26'd13731; ROM2[72]<=26'd17917; ROM3[72]<=26'd32347; ROM4[72]<=26'd18083;
ROM1[73]<=26'd15482; ROM2[73]<=26'd17535; ROM3[73]<=26'd29215; ROM4[73]<=26'd32781;
ROM1[74]<=-26'd3839; ROM2[74]<=-26'd2363; ROM3[74]<=26'd5655; ROM4[74]<=-26'd21117;
ROM1[75]<=26'd45895; ROM2[75]<=26'd54021; ROM3[75]<=26'd70162; ROM4[75]<=26'd99153;
ROM1[76]<=26'd61012; ROM2[76]<=26'd68377; ROM3[76]<=26'd87495; ROM4[76]<=26'd145944;
ROM1[77]<=26'd8874; ROM2[77]<=26'd12210; ROM3[77]<=26'd25858; ROM4[77]<=26'd7438;
ROM1[78]<=26'd23571; ROM2[78]<=26'd30856; ROM3[78]<=26'd51399; ROM4[78]<=26'd33339;
ROM1[79]<=26'd18019; ROM2[79]<=26'd22682; ROM3[79]<=26'd44225; ROM4[79]<=26'd26080;
ROM1[80]<=26'd23500; ROM2[80]<=26'd27114; ROM3[80]<=26'd53205; ROM4[80]<=26'd44244;
ROM1[81]<=26'd22242; ROM2[81]<=26'd28300; ROM3[81]<=26'd55605; ROM4[81]<=26'd30750;
ROM1[82]<=26'd21062; ROM2[82]<=26'd26141; ROM3[82]<=26'd51747; ROM4[82]<=26'd31775;
ROM1[83]<=26'd17775; ROM2[83]<=26'd21911; ROM3[83]<=26'd44183; ROM4[83]<=26'd27155;
ROM1[84]<=26'd16917; ROM2[84]<=26'd23971; ROM3[84]<=26'd50298; ROM4[84]<=26'd11651;
ROM1[85]<=26'd21705; ROM2[85]<=26'd27147; ROM3[85]<=26'd58810; ROM4[85]<=26'd29412;
ROM1[86]<=26'd19288; ROM2[86]<=26'd24208; ROM3[86]<=26'd53200; ROM4[86]<=26'd25469;
ROM1[87]<=26'd17835; ROM2[87]<=26'd23329; ROM3[87]<=26'd50557; ROM4[87]<=26'd19852;
ROM1[88]<=26'd16523; ROM2[88]<=26'd21782; ROM3[88]<=26'd49990; ROM4[88]<=26'd16300;
ROM1[89]<=26'd9698; ROM2[89]<=26'd16475; ROM3[89]<=26'd43768; ROM4[89]<=-26'd9422;
ROM1[90]<=26'd15346; ROM2[90]<=26'd23219; ROM3[90]<=26'd57110; ROM4[90]<=26'd97;
ROM1[91]<=26'd16963; ROM2[91]<=26'd24746; ROM3[91]<=26'd60102; ROM4[91]<=26'd4526;
ROM1[92]<=26'd16228; ROM2[92]<=26'd24029; ROM3[92]<=26'd62668; ROM4[92]<=26'd576;
ROM1[93]<=26'd20079; ROM2[93]<=26'd30732; ROM3[93]<=26'd75232; ROM4[93]<=-26'd1537;
ROM1[94]<=26'd26946; ROM2[94]<=26'd35178; ROM3[94]<=26'd81357; ROM4[94]<=26'd27248;
ROM1[95]<=26'd19540; ROM2[95]<=26'd24193; ROM3[95]<=26'd69310; ROM4[95]<=26'd18926;
ROM1[96]<=26'd30123; ROM2[96]<=26'd36163; ROM3[96]<=26'd84082; ROM4[96]<=26'd44015;
ROM1[97]<=26'd6811; ROM2[97]<=26'd9042; ROM3[97]<=26'd54397; ROM4[97]<=-26'd10421;
ROM1[98]<=26'd127176; ROM2[98]<=26'd144399; ROM3[98]<=26'd217318; ROM4[98]<=26'd280602;
ROM1[99]<=26'd131912; ROM2[99]<=26'd151404; ROM3[99]<=26'd228097; ROM4[99]<=26'd284344;
ROM1[100]<=26'd36432; ROM2[100]<=26'd44964; ROM3[100]<=26'd101753; ROM4[100]<=26'd48890;
ROM1[101]<=26'd38079; ROM2[101]<=26'd44472; ROM3[101]<=26'd102580; ROM4[101]<=26'd61120;
ROM1[102]<=26'd22281; ROM2[102]<=26'd24700; ROM3[102]<=26'd81684; ROM4[102]<=26'd29122;
ROM1[103]<=26'd43720; ROM2[103]<=26'd51824; ROM3[103]<=26'd115446; ROM4[103]<=26'd68734;
ROM1[104]<=26'd36464; ROM2[104]<=26'd44758; ROM3[104]<=26'd110315; ROM4[104]<=26'd45227;
ROM1[105]<=26'd37596; ROM2[105]<=26'd46034; ROM3[105]<=26'd113752; ROM4[105]<=26'd46946;
ROM1[106]<=26'd48706; ROM2[106]<=26'd60458; ROM3[106]<=26'd134293; ROM4[106]<=26'd64731;
ROM1[107]<=26'd39269; ROM2[107]<=26'd46853; ROM3[107]<=26'd116445; ROM4[107]<=26'd54131;
ROM1[108]<=26'd31897; ROM2[108]<=26'd37263; ROM3[108]<=26'd104138; ROM4[108]<=26'd41651;
ROM1[109]<=26'd24172; ROM2[109]<=26'd24810; ROM3[109]<=26'd86214; ROM4[109]<=26'd38905;
ROM1[110]<=26'd26060; ROM2[110]<=26'd27203; ROM3[110]<=26'd90735; ROM4[110]<=26'd41591;
ROM1[111]<=26'd39041; ROM2[111]<=26'd42771; ROM3[111]<=26'd111789; ROM4[111]<=26'd68074;
ROM1[112]<=26'd41505; ROM2[112]<=26'd46783; ROM3[112]<=26'd116085; ROM4[112]<=26'd69509;
ROM1[113]<=26'd42734; ROM2[113]<=26'd52007; ROM3[113]<=26'd123943; ROM4[113]<=26'd56906;
ROM1[114]<=26'd36083; ROM2[114]<=26'd39532; ROM3[114]<=26'd107101; ROM4[114]<=26'd60982;
ROM1[115]<=26'd41492; ROM2[115]<=26'd48970; ROM3[115]<=26'd119467; ROM4[115]<=26'd60657;
ROM1[116]<=26'd32705; ROM2[116]<=26'd38570; ROM3[116]<=26'd107114; ROM4[116]<=26'd41351;
ROM1[117]<=26'd39777; ROM2[117]<=26'd45222; ROM3[117]<=26'd118654; ROM4[117]<=26'd61731;
ROM1[118]<=26'd44696; ROM2[118]<=26'd53497; ROM3[118]<=26'd128405; ROM4[118]<=26'd63213;
ROM1[119]<=26'd43144; ROM2[119]<=26'd52521; ROM3[119]<=26'd126328; ROM4[119]<=26'd56999;
ROM1[120]<=26'd47882; ROM2[120]<=26'd57709; ROM3[120]<=26'd134435; ROM4[120]<=26'd68123;
ROM1[121]<=26'd46692; ROM2[121]<=26'd56817; ROM3[121]<=26'd135354; ROM4[121]<=26'd62587;
ROM1[122]<=26'd54617; ROM2[122]<=26'd68871; ROM3[122]<=26'd151086; ROM4[122]<=26'd69105;
ROM1[123]<=26'd64578; ROM2[123]<=26'd83434; ROM3[123]<=26'd173301; ROM4[123]<=26'd77974;
ROM1[124]<=26'd67714; ROM2[124]<=26'd89350; ROM3[124]<=26'd181821; ROM4[124]<=26'd75726;
ROM1[125]<=26'd67909; ROM2[125]<=26'd87820; ROM3[125]<=26'd174664; ROM4[125]<=26'd85665;
ROM1[126]<=26'd59091; ROM2[126]<=26'd76750; ROM3[126]<=26'd154043; ROM4[126]<=26'd72499;
ROM1[127]<=26'd67239; ROM2[127]<=26'd89551; ROM3[127]<=26'd176634; ROM4[127]<=26'd74663;



/*
        ROM1[0]<=-26'd3696; ROM2[0]<=-26'd11888; ROM3[0]<=26'd800; ROM4[0]<=26'd8603;
        ROM1[1]<=26'd7920; ROM2[1]<=-26'd2203; ROM3[1]<=26'd17669; ROM4[1]<=26'd42064;
        ROM1[2]<=26'd9044; ROM2[2]<=26'd1067; ROM3[2]<=26'd17670; ROM4[2]<=26'd41552;
        ROM1[3]<=26'd10583; ROM2[3]<=26'd4716; ROM3[3]<=26'd18538; ROM4[3]<=26'd42808;
        ROM1[4]<=26'd11555; ROM2[4]<=26'd7746; ROM3[4]<=26'd18330; ROM4[4]<=26'd41840;
        ROM1[5]<=26'd15277; ROM2[5]<=26'd13458; ROM3[5]<=26'd23699; ROM4[5]<=26'd52283;
        ROM1[6]<=26'd15396; ROM2[6]<=26'd15482; ROM3[6]<=26'd21953; ROM4[6]<=26'd48112;
        ROM1[7]<=26'd20854; ROM2[7]<=26'd22746; ROM3[7]<=26'd30990; ROM4[7]<=26'd66015;
        ROM1[8]<=26'd23079; ROM2[8]<=26'd26668; ROM3[8]<=26'd33684; ROM4[8]<=26'd70876;
        ROM1[9]<=26'd19852; ROM2[9]<=26'd25017; ROM3[9]<=26'd25605; ROM4[9]<=26'd53615;
        ROM1[10]<=26'd24606; ROM2[10]<=26'd31217; ROM3[10]<=26'd33628; ROM4[10]<=26'd69320;
        ROM1[11]<=26'd23738; ROM2[11]<=26'd31660; ROM3[11]<=26'd30556; ROM4[11]<=26'd62237;
        ROM1[12]<=26'd25216; ROM2[12]<=26'd34308; ROM3[12]<=26'd32330; ROM4[12]<=26'd65042;
        ROM1[13]<=26'd29173; ROM2[13]<=26'd39293; ROM3[13]<=26'd39217; ROM4[13]<=26'd78281;
        ROM1[14]<=26'd23071; ROM2[14]<=26'd34076; ROM3[14]<=26'd26141; ROM4[14]<=26'd50550;
        ROM1[15]<=26'd23974; ROM2[15]<=26'd35723; ROM3[15]<=26'd27228; ROM4[15]<=26'd51807;
        ROM1[16]<=26'd7689; ROM2[16]<=26'd3664; ROM3[16]<=26'd10472; ROM4[16]<=26'd30368;
        ROM1[17]<=-26'd1509; ROM2[17]<=26'd3138; ROM3[17]<=-26'd163; ROM4[17]<=26'd8738;
        ROM1[18]<=-26'd1534; ROM2[18]<=26'd3473; ROM3[18]<=-26'd512; ROM4[18]<=26'd6925;
        ROM1[19]<=-26'd460; ROM2[19]<=26'd4797; ROM3[19]<=26'd1457; ROM4[19]<=26'd9828;
        ROM1[20]<=26'd663; ROM2[20]<=26'd6074; ROM3[20]<=26'd3629; ROM4[20]<=26'd13116;
        ROM1[21]<=-26'd650; ROM2[21]<=26'd4831; ROM3[21]<=26'd1021; ROM4[21]<=26'd6579;
        ROM1[22]<=-26'd3320; ROM2[22]<=26'd2163; ROM3[22]<=-26'd4228; ROM4[22]<=-26'd5397;
        ROM1[23]<=-26'd658; ROM2[23]<=26'd4776; ROM3[23]<=26'd1245; ROM4[23]<=26'd4591;
        ROM1[24]<=-26'd6065; ROM2[24]<=-26'd715; ROM3[24]<=-26'd9385; ROM4[24]<=-26'd18443;
        ROM1[25]<=-26'd1790; ROM2[25]<=26'd3460; ROM3[25]<=-26'd630; ROM4[25]<=-26'd1743;
        ROM1[26]<=-26'd5854; ROM2[26]<=-26'd705; ROM3[26]<=-26'd8557; ROM4[26]<=-26'd19241;
        ROM1[27]<=26'd731; ROM2[27]<=26'd5800; ROM3[27]<=26'd4794; ROM4[27]<=26'd6889;
        ROM1[28]<=-26'd2679; ROM2[28]<=26'd2346; ROM3[28]<=-26'd1883; ROM4[28]<=-26'd8030;
        ROM1[29]<=-26'd3454; ROM2[29]<=26'd1581; ROM3[29]<=-26'd3351; ROM4[29]<=-26'd12250;
        ROM1[30]<=-26'd4518; ROM2[30]<=26'd598; ROM3[30]<=-26'd5471; ROM4[30]<=-26'd17785;
        ROM1[31]<=-26'd98; ROM2[31]<=26'd5182; ROM3[31]<=26'd3282; ROM4[31]<=-26'd1004;
        ROM1[32]<=-26'd18754; ROM2[32]<=-26'd29594; ROM3[32]<=-26'd17841; ROM4[32]<=-26'd31507;
        ROM1[33]<=-26'd17400; ROM2[33]<=-26'd27865; ROM3[33]<=-26'd15447; ROM4[33]<=-26'd27692;
        ROM1[34]<=-26'd4974; ROM2[34]<=-26'd23135; ROM3[34]<=26'd766; ROM4[34]<=26'd3263;
        ROM1[35]<=26'd595; ROM2[35]<=-26'd16940; ROM3[35]<=26'd11314; ROM4[35]<=26'd23877;
        ROM1[36]<=26'd1336; ROM2[36]<=-26'd15436; ROM3[36]<=26'd12060; ROM4[36]<=26'd24440;
        ROM1[37]<=26'd2291; ROM2[37]<=-26'd13578; ROM3[37]<=26'd13077; ROM4[37]<=26'd25606;
        ROM1[38]<=26'd6013; ROM2[38]<=-26'd8811; ROM3[38]<=26'd19474; ROM4[38]<=26'd37846;
        ROM1[39]<=26'd5041; ROM2[39]<=-26'd8594; ROM3[39]<=26'd16328; ROM4[39]<=26'd30571;
        ROM1[40]<=26'd3702; ROM2[40]<=-26'd8606; ROM3[40]<=26'd12294; ROM4[40]<=26'd21522;
        ROM1[41]<=26'd5761; ROM2[41]<=-26'd5083; ROM3[41]<=26'd14910; ROM4[41]<=26'd26148;
        ROM1[42]<=26'd9437; ROM2[42]<=26'd185; ROM3[42]<=26'd20619; ROM4[42]<=26'd37157;
        ROM1[43]<=26'd5865; ROM2[43]<=-26'd1676; ROM3[43]<=26'd11702; ROM4[43]<=26'd18222;
        ROM1[44]<=26'd12582; ROM2[44]<=26'd6861; ROM3[44]<=26'd23245; ROM4[44]<=26'd41266;
        ROM1[45]<=26'd14450; ROM2[45]<=26'd10646; ROM3[45]<=26'd24983; ROM4[45]<=26'd44242;
        ROM1[46]<=26'd12590; ROM2[46]<=26'd10785; ROM3[46]<=26'd19178; ROM4[46]<=26'd31780;
        ROM1[47]<=26'd13895; ROM2[47]<=26'd14155; ROM3[47]<=26'd19627; ROM4[47]<=26'd32161;
        ROM1[48]<=26'd1056; ROM2[48]<=-26'd12951; ROM3[48]<=26'd8119; ROM4[48]<=26'd21974;
        ROM1[49]<=26'd3500; ROM2[49]<=-26'd8358; ROM3[49]<=26'd10755; ROM4[49]<=26'd26867;
        ROM1[50]<=-26'd9131; ROM2[50]<=-26'd10631; ROM3[50]<=-26'd8582; ROM4[50]<=-26'd12051;
        ROM1[51]<=-26'd8148; ROM2[51]<=-26'd7486; ROM3[51]<=-26'd8883; ROM4[51]<=-26'd13176;
        ROM1[52]<=-26'd1603; ROM2[52]<=26'd1203; ROM3[52]<=26'd1964; ROM4[52]<=26'd8547;
        ROM1[53]<=-26'd6856; ROM2[53]<=-26'd1946; ROM3[53]<=-26'd10745; ROM4[53]<=-26'd18033;
        ROM1[54]<=-26'd4023; ROM2[54]<=26'd2937; ROM3[54]<=-26'd7222; ROM4[54]<=-26'd11355;
        ROM1[55]<=-26'd2520; ROM2[55]<=26'd6420; ROM3[55]<=-26'd6281; ROM4[55]<=-26'd9992;
        ROM1[56]<=26'd3324; ROM2[56]<=26'd14157; ROM3[56]<=26'd3435; ROM4[56]<=26'd9330;
        ROM1[57]<=26'd1773; ROM2[57]<=26'd14400; ROM3[57]<=-26'd1529; ROM4[57]<=-26'd1476;
        ROM1[58]<=26'd5141; ROM2[58]<=26'd19449; ROM3[58]<=26'd3465; ROM4[58]<=26'd8099;
        ROM1[59]<=26'd4835; ROM2[59]<=26'd20703; ROM3[59]<=26'd1246; ROM4[59]<=26'd2845;
        ROM1[60]<=26'd5528; ROM2[60]<=26'd22826; ROM3[60]<=26'd1167; ROM4[60]<=26'd1936;
        ROM1[61]<=26'd6399; ROM2[61]<=26'd24990; ROM3[61]<=26'd1593; ROM4[61]<=26'd2016;
        ROM1[62]<=26'd12013; ROM2[62]<=26'd31756; ROM3[62]<=26'd11657; ROM4[62]<=26'd21810;
        ROM1[63]<=26'd8780; ROM2[63]<=26'd29532; ROM3[63]<=26'd4183; ROM4[63]<=26'd5604;
        ROM1[64]<=-26'd6244; ROM2[64]<=-26'd1009; ROM3[64]<=-26'd10332; ROM4[64]<=-26'd11157;
        ROM1[65]<=-26'd4079; ROM2[65]<=26'd1884; ROM3[65]<=-26'd6701; ROM4[65]<=-26'd4691;
        ROM1[66]<=26'd259; ROM2[66]<=26'd6813; ROM3[66]<=26'd1421; ROM4[66]<=26'd10938;
        ROM1[67]<=26'd11229; ROM2[67]<=26'd10056; ROM3[67]<=26'd14756; ROM4[67]<=26'd35983;
        ROM1[68]<=26'd17705; ROM2[68]<=26'd16878; ROM3[68]<=26'd27427; ROM4[68]<=26'd60856;
        ROM1[69]<=26'd11938; ROM2[69]<=26'd11348; ROM3[69]<=26'd15726; ROM4[69]<=26'd35734;
        ROM1[70]<=26'd19373; ROM2[70]<=26'd18925; ROM3[70]<=26'd30535; ROM4[70]<=26'd64923;
        ROM1[71]<=26'd15362; ROM2[71]<=26'd14975; ROM3[71]<=26'd22541; ROM4[71]<=26'd47339;
        ROM1[72]<=26'd19613; ROM2[72]<=26'd19221; ROM3[72]<=26'd31143; ROM4[72]<=26'd63758;
        ROM1[73]<=26'd16611; ROM2[73]<=26'd16163; ROM3[73]<=26'd25291; ROM4[73]<=26'd50528;
        ROM1[74]<=26'd17726; ROM2[74]<=26'd17192; ROM3[74]<=26'd27712; ROM4[74]<=26'd54247;
        ROM1[75]<=26'd11993; ROM2[75]<=26'd11357; ROM3[75]<=26'd16449; ROM4[75]<=26'd29910;
        ROM1[76]<=26'd13993; ROM2[76]<=26'd13259; ROM3[76]<=26'd20651; ROM4[76]<=26'd37276;
        ROM1[77]<=26'd12685; ROM2[77]<=26'd11874; ROM3[77]<=26'd18212; ROM4[77]<=26'd31037;
        ROM1[78]<=26'd14186; ROM2[78]<=26'd13337; ROM3[78]<=26'd21349; ROM4[78]<=26'd36240;
        ROM1[79]<=26'd12843; ROM2[79]<=26'd12012; ROM3[79]<=26'd18737; ROM4[79]<=26'd29676;
        ROM1[80]<=-26'd1734; ROM2[80]<=-26'd18858; ROM3[80]<=26'd5964; ROM4[80]<=26'd16233;
        ROM1[81]<=-26'd690; ROM2[81]<=-26'd17638; ROM3[81]<=26'd7952; ROM4[81]<=26'd19150;
        ROM1[82]<=-26'd3212; ROM2[82]<=-26'd19883; ROM3[82]<=26'd2698; ROM4[82]<=26'd7257;
        ROM1[83]<=26'd2383; ROM2[83]<=-26'd13898; ROM3[83]<=26'd13558; ROM4[83]<=26'd28431;
        ROM1[84]<=-26'd14473; ROM2[84]<=-26'd22049; ROM3[84]<=-26'd12426; ROM4[84]<=-26'd24655;
        ROM1[85]<=-26'd16262; ROM2[85]<=-26'd23195; ROM3[85]<=-26'd16612; ROM4[85]<=-26'd34241;
        ROM1[86]<=-26'd13346; ROM2[86]<=-26'd19500; ROM3[86]<=-26'd11539; ROM4[86]<=-26'd24799;
        ROM1[87]<=-26'd15932; ROM2[87]<=-26'd21164; ROM3[87]<=-26'd17621; ROM4[87]<=-26'd38182;
        ROM1[88]<=-26'd10922; ROM2[88]<=-26'd15091; ROM3[88]<=-26'd8669; ROM4[88]<=-26'd20696;
        ROM1[89]<=-26'd6837; ROM2[89]<=-26'd9800; ROM3[89]<=-26'd1721; ROM4[89]<=-26'd7273;
        ROM1[90]<=-26'd10523; ROM2[90]<=-26'd12140; ROM3[90]<=-26'd10467; ROM4[90]<=-26'd25977;
        ROM1[91]<=-26'd6226; ROM2[91]<=-26'd6363; ROM3[91]<=-26'd3393; ROM4[91]<=-26'd12208;
        ROM1[92]<=-26'd9059; ROM2[92]<=-26'd7588; ROM3[92]<=-26'd10718; ROM4[92]<=-26'd27913;
        ROM1[93]<=-26'd2608; ROM2[93]<=26'd589; ROM3[93]<=26'd395; ROM4[93]<=-26'd5780;
        ROM1[94]<=-26'd4345; ROM2[94]<=26'd685; ROM3[94]<=-26'd4985; ROM4[94]<=-26'd17424;
        ROM1[95]<=-26'd3368; ROM2[95]<=26'd3589; ROM3[95]<=-26'd5042; ROM4[95]<=-26'd18125;
        ROM1[96]<=-26'd14529; ROM2[96]<=-26'd21947; ROM3[96]<=-26'd13076; ROM4[96]<=-26'd21226;
        ROM1[97]<=-26'd17191; ROM2[97]<=-26'd22536; ROM3[97]<=-26'd20566; ROM4[97]<=-26'd37119;
        ROM1[98]<=-26'd8542; ROM2[98]<=-26'd11766; ROM3[98]<=-26'd5490; ROM4[98]<=-26'd6733;
        ROM1[99]<=-26'd13244; ROM2[99]<=-26'd14315; ROM3[99]<=-26'd17148; ROM4[99]<=-26'd31141;
        ROM1[100]<=26'd10718; ROM2[100]<=26'd3621; ROM3[100]<=26'd20314; ROM4[100]<=26'd43919;
        ROM1[101]<=26'd9436; ROM2[101]<=26'd4500; ROM3[101]<=26'd15486; ROM4[101]<=26'd33514;
        ROM1[102]<=26'd15285; ROM2[102]<=26'd12488; ROM3[102]<=26'd24944; ROM4[102]<=26'd52390;
        ROM1[103]<=26'd19146; ROM2[103]<=26'd18449; ROM3[103]<=26'd30471; ROM4[103]<=26'd63192;
        ROM1[104]<=26'd15252; ROM2[104]<=26'd16596; ROM3[104]<=26'd20549; ROM4[104]<=26'd42304;
        ROM1[105]<=26'd19818; ROM2[105]<=26'd23132; ROM3[105]<=26'd27627; ROM4[105]<=26'd56243;
        ROM1[106]<=26'd21752; ROM2[106]<=26'd26947; ROM3[106]<=26'd29537; ROM4[106]<=26'd59559;
        ROM1[107]<=26'd23302; ROM2[107]<=26'd30277; ROM3[107]<=26'd30788; ROM4[107]<=26'd61493;
        ROM1[108]<=26'd22051; ROM2[108]<=26'd30693; ROM3[108]<=26'd26561; ROM4[108]<=26'd52158;
        ROM1[109]<=26'd29525; ROM2[109]<=26'd39711; ROM3[109]<=26'd39920; ROM4[109]<=26'd78834;
        ROM1[110]<=26'd26761; ROM2[110]<=26'd38359; ROM3[110]<=26'd32945; ROM4[110]<=26'd63782;
        ROM1[111]<=26'd31285; ROM2[111]<=26'd44158; ROM3[111]<=26'd40696; ROM4[111]<=26'd78873;
        ROM1[112]<=26'd14822; ROM2[112]<=26'd12445; ROM3[112]<=26'd23011; ROM4[112]<=26'd55701;
        ROM1[113]<=26'd12524; ROM2[113]<=26'd11138; ROM3[113]<=26'd17426; ROM4[113]<=26'd43362;
        ROM1[114]<=26'd17619; ROM2[114]<=26'd17082; ROM3[114]<=26'd26785; ROM4[114]<=26'd61610;
        ROM1[115]<=26'd14940; ROM2[115]<=26'd15113; ROM3[115]<=26'd20746; ROM4[115]<=26'd48247;
        ROM1[116]<=26'd19527; ROM2[116]<=26'd20275; ROM3[116]<=26'd29385; ROM4[116]<=26'd64932;
        ROM1[117]<=26'd1188; ROM2[117]<=26'd10578; ROM3[117]<=26'd505; ROM4[117]<=26'd5888;
        ROM1[118]<=26'd4045; ROM2[118]<=26'd13765; ROM3[118]<=26'd5950; ROM4[118]<=26'd15943;
        ROM1[119]<=26'd2793; ROM2[119]<=26'd12738; ROM3[119]<=26'd3295; ROM4[119]<=26'd9359;
        ROM1[120]<=26'd3274; ROM2[120]<=26'd13349; ROM3[120]<=26'd4207; ROM4[120]<=26'd10058;
        ROM1[121]<=26'd1580; ROM2[121]<=26'd11707; ROM3[121]<=26'd857; ROM4[121]<=26'd1992;
        ROM1[122]<=26'd5388; ROM2[122]<=26'd15502; ROM3[122]<=26'd8581; ROM4[122]<=26'd16605;
        ROM1[123]<=26'd2870; ROM2[123]<=26'd12925; ROM3[123]<=26'd3705; ROM4[123]<=26'd5376;
        ROM1[124]<=26'd1079; ROM2[124]<=26'd11044; ROM3[124]<=26'd315; ROM4[124]<=-26'd2819;
        ROM1[125]<=26'd2575; ROM2[125]<=26'd12438; ROM3[125]<=26'd3513; ROM4[125]<=26'd2488;
        ROM1[126]<=-26'd2229; ROM2[126]<=26'd7538; ROM3[126]<=-26'd5897; ROM4[126]<=-26'd18048;
        ROM1[127]<=-26'd16272; ROM2[127]<=-26'd22962; ROM3[127]<=-26'd17426; ROM4[127]<=-26'd28994;
*/


	end
	else begin
		if(cnt == 7'd127) begin
				cnt<=0;
			end
		//?��?��?�� addr?��?��.
		data1 <= ROM1[cnt];
		data2 <= ROM2[cnt];
		data3 <= ROM3[cnt];
		data4 <= ROM4[cnt];
		cnt <= cnt+1'b1;
	end
end
endmodule 
