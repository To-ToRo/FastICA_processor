//출처 : https://verilogguide.readthedocs.io/en/latest/verilog/designs.html#read-only-memory-rom

module ROM(
    input wire clk,
	input wire En,
    input wire  [13:0] addr,
    output reg signed [25:0] data1,
	output reg signed [25:0] data2,
	output reg signed [25:0] data3,
	output reg signed [25:0] data4
);

//ROM[0]?�� ?���? : 16bit(?�� ?��그널?�� ?���?) * 4(4개의 ?��그널) 
// 각각?�� ?��그널?�� �? 1000sample?�� ?��?���?�? addr??  16비트�? ?��?��(0~39999 < 0~65536) 

reg signed [25:0] ROM1[0:127];
reg signed [25:0] ROM2[0:127];
reg signed [25:0] ROM3[0:127];
reg signed [25:0] ROM4[0:127];
reg [6:0] cnt;

always @(posedge clk) begin
	if(!En) begin
		cnt<=0;
        data1<=0;
        data2<=0;
        data3<=0;
        data4<=0;

        ROM1[0]<=-26'd3696; ROM2[0]<=-26'd11888; ROM3[0]<=26'd800; ROM4[0]<=26'd8603;
        ROM1[1]<=26'd7920; ROM2[1]<=-26'd2203; ROM3[1]<=26'd17669; ROM4[1]<=26'd42064;
        ROM1[2]<=26'd9044; ROM2[2]<=26'd1067; ROM3[2]<=26'd17670; ROM4[2]<=26'd41552;
        ROM1[3]<=26'd10583; ROM2[3]<=26'd4716; ROM3[3]<=26'd18538; ROM4[3]<=26'd42808;
        ROM1[4]<=26'd11555; ROM2[4]<=26'd7746; ROM3[4]<=26'd18330; ROM4[4]<=26'd41840;
        ROM1[5]<=26'd15277; ROM2[5]<=26'd13458; ROM3[5]<=26'd23699; ROM4[5]<=26'd52283;
        ROM1[6]<=26'd15396; ROM2[6]<=26'd15482; ROM3[6]<=26'd21953; ROM4[6]<=26'd48112;
        ROM1[7]<=26'd20854; ROM2[7]<=26'd22746; ROM3[7]<=26'd30990; ROM4[7]<=26'd66015;
        ROM1[8]<=26'd23079; ROM2[8]<=26'd26668; ROM3[8]<=26'd33684; ROM4[8]<=26'd70876;
        ROM1[9]<=26'd19852; ROM2[9]<=26'd25017; ROM3[9]<=26'd25605; ROM4[9]<=26'd53615;
        ROM1[10]<=26'd24606; ROM2[10]<=26'd31217; ROM3[10]<=26'd33628; ROM4[10]<=26'd69320;
        ROM1[11]<=26'd23738; ROM2[11]<=26'd31660; ROM3[11]<=26'd30556; ROM4[11]<=26'd62237;
        ROM1[12]<=26'd25216; ROM2[12]<=26'd34308; ROM3[12]<=26'd32330; ROM4[12]<=26'd65042;
        ROM1[13]<=26'd29173; ROM2[13]<=26'd39293; ROM3[13]<=26'd39217; ROM4[13]<=26'd78281;
        ROM1[14]<=26'd23071; ROM2[14]<=26'd34076; ROM3[14]<=26'd26141; ROM4[14]<=26'd50550;
        ROM1[15]<=26'd23974; ROM2[15]<=26'd35723; ROM3[15]<=26'd27228; ROM4[15]<=26'd51807;
        ROM1[16]<=26'd7689; ROM2[16]<=26'd3664; ROM3[16]<=26'd10472; ROM4[16]<=26'd30368;
        ROM1[17]<=-26'd1509; ROM2[17]<=26'd3138; ROM3[17]<=-26'd163; ROM4[17]<=26'd8738;
        ROM1[18]<=-26'd1534; ROM2[18]<=26'd3473; ROM3[18]<=-26'd512; ROM4[18]<=26'd6925;
        ROM1[19]<=-26'd460; ROM2[19]<=26'd4797; ROM3[19]<=26'd1457; ROM4[19]<=26'd9828;
        ROM1[20]<=26'd663; ROM2[20]<=26'd6074; ROM3[20]<=26'd3629; ROM4[20]<=26'd13116;
        ROM1[21]<=-26'd650; ROM2[21]<=26'd4831; ROM3[21]<=26'd1021; ROM4[21]<=26'd6579;
        ROM1[22]<=-26'd3320; ROM2[22]<=26'd2163; ROM3[22]<=-26'd4228; ROM4[22]<=-26'd5397;
        ROM1[23]<=-26'd658; ROM2[23]<=26'd4776; ROM3[23]<=26'd1245; ROM4[23]<=26'd4591;
        ROM1[24]<=-26'd6065; ROM2[24]<=-26'd715; ROM3[24]<=-26'd9385; ROM4[24]<=-26'd18443;
        ROM1[25]<=-26'd1790; ROM2[25]<=26'd3460; ROM3[25]<=-26'd630; ROM4[25]<=-26'd1743;
        ROM1[26]<=-26'd5854; ROM2[26]<=-26'd705; ROM3[26]<=-26'd8557; ROM4[26]<=-26'd19241;
        ROM1[27]<=26'd731; ROM2[27]<=26'd5800; ROM3[27]<=26'd4794; ROM4[27]<=26'd6889;
        ROM1[28]<=-26'd2679; ROM2[28]<=26'd2346; ROM3[28]<=-26'd1883; ROM4[28]<=-26'd8030;
        ROM1[29]<=-26'd3454; ROM2[29]<=26'd1581; ROM3[29]<=-26'd3351; ROM4[29]<=-26'd12250;
        ROM1[30]<=-26'd4518; ROM2[30]<=26'd598; ROM3[30]<=-26'd5471; ROM4[30]<=-26'd17785;
        ROM1[31]<=-26'd98; ROM2[31]<=26'd5182; ROM3[31]<=26'd3282; ROM4[31]<=-26'd1004;
        ROM1[32]<=-26'd18754; ROM2[32]<=-26'd29594; ROM3[32]<=-26'd17841; ROM4[32]<=-26'd31507;
        ROM1[33]<=-26'd17400; ROM2[33]<=-26'd27865; ROM3[33]<=-26'd15447; ROM4[33]<=-26'd27692;
        ROM1[34]<=-26'd4974; ROM2[34]<=-26'd23135; ROM3[34]<=26'd766; ROM4[34]<=26'd3263;
        ROM1[35]<=26'd595; ROM2[35]<=-26'd16940; ROM3[35]<=26'd11314; ROM4[35]<=26'd23877;
        ROM1[36]<=26'd1336; ROM2[36]<=-26'd15436; ROM3[36]<=26'd12060; ROM4[36]<=26'd24440;
        ROM1[37]<=26'd2291; ROM2[37]<=-26'd13578; ROM3[37]<=26'd13077; ROM4[37]<=26'd25606;
        ROM1[38]<=26'd6013; ROM2[38]<=-26'd8811; ROM3[38]<=26'd19474; ROM4[38]<=26'd37846;
        ROM1[39]<=26'd5041; ROM2[39]<=-26'd8594; ROM3[39]<=26'd16328; ROM4[39]<=26'd30571;
        ROM1[40]<=26'd3702; ROM2[40]<=-26'd8606; ROM3[40]<=26'd12294; ROM4[40]<=26'd21522;
        ROM1[41]<=26'd5761; ROM2[41]<=-26'd5083; ROM3[41]<=26'd14910; ROM4[41]<=26'd26148;
        ROM1[42]<=26'd9437; ROM2[42]<=26'd185; ROM3[42]<=26'd20619; ROM4[42]<=26'd37157;
        ROM1[43]<=26'd5865; ROM2[43]<=-26'd1676; ROM3[43]<=26'd11702; ROM4[43]<=26'd18222;
        ROM1[44]<=26'd12582; ROM2[44]<=26'd6861; ROM3[44]<=26'd23245; ROM4[44]<=26'd41266;
        ROM1[45]<=26'd14450; ROM2[45]<=26'd10646; ROM3[45]<=26'd24983; ROM4[45]<=26'd44242;
        ROM1[46]<=26'd12590; ROM2[46]<=26'd10785; ROM3[46]<=26'd19178; ROM4[46]<=26'd31780;
        ROM1[47]<=26'd13895; ROM2[47]<=26'd14155; ROM3[47]<=26'd19627; ROM4[47]<=26'd32161;
        ROM1[48]<=26'd1056; ROM2[48]<=-26'd12951; ROM3[48]<=26'd8119; ROM4[48]<=26'd21974;
        ROM1[49]<=26'd3500; ROM2[49]<=-26'd8358; ROM3[49]<=26'd10755; ROM4[49]<=26'd26867;
        ROM1[50]<=-26'd9131; ROM2[50]<=-26'd10631; ROM3[50]<=-26'd8582; ROM4[50]<=-26'd12051;
        ROM1[51]<=-26'd8148; ROM2[51]<=-26'd7486; ROM3[51]<=-26'd8883; ROM4[51]<=-26'd13176;
        ROM1[52]<=-26'd1603; ROM2[52]<=26'd1203; ROM3[52]<=26'd1964; ROM4[52]<=26'd8547;
        ROM1[53]<=-26'd6856; ROM2[53]<=-26'd1946; ROM3[53]<=-26'd10745; ROM4[53]<=-26'd18033;
        ROM1[54]<=-26'd4023; ROM2[54]<=26'd2937; ROM3[54]<=-26'd7222; ROM4[54]<=-26'd11355;
        ROM1[55]<=-26'd2520; ROM2[55]<=26'd6420; ROM3[55]<=-26'd6281; ROM4[55]<=-26'd9992;
        ROM1[56]<=26'd3324; ROM2[56]<=26'd14157; ROM3[56]<=26'd3435; ROM4[56]<=26'd9330;
        ROM1[57]<=26'd1773; ROM2[57]<=26'd14400; ROM3[57]<=-26'd1529; ROM4[57]<=-26'd1476;
        ROM1[58]<=26'd5141; ROM2[58]<=26'd19449; ROM3[58]<=26'd3465; ROM4[58]<=26'd8099;
        ROM1[59]<=26'd4835; ROM2[59]<=26'd20703; ROM3[59]<=26'd1246; ROM4[59]<=26'd2845;
        ROM1[60]<=26'd5528; ROM2[60]<=26'd22826; ROM3[60]<=26'd1167; ROM4[60]<=26'd1936;
        ROM1[61]<=26'd6399; ROM2[61]<=26'd24990; ROM3[61]<=26'd1593; ROM4[61]<=26'd2016;
        ROM1[62]<=26'd12013; ROM2[62]<=26'd31756; ROM3[62]<=26'd11657; ROM4[62]<=26'd21810;
        ROM1[63]<=26'd8780; ROM2[63]<=26'd29532; ROM3[63]<=26'd4183; ROM4[63]<=26'd5604;
        ROM1[64]<=-26'd6244; ROM2[64]<=-26'd1009; ROM3[64]<=-26'd10332; ROM4[64]<=-26'd11157;
        ROM1[65]<=-26'd4079; ROM2[65]<=26'd1884; ROM3[65]<=-26'd6701; ROM4[65]<=-26'd4691;
        ROM1[66]<=26'd259; ROM2[66]<=26'd6813; ROM3[66]<=26'd1421; ROM4[66]<=26'd10938;
        ROM1[67]<=26'd11229; ROM2[67]<=26'd10056; ROM3[67]<=26'd14756; ROM4[67]<=26'd35983;
        ROM1[68]<=26'd17705; ROM2[68]<=26'd16878; ROM3[68]<=26'd27427; ROM4[68]<=26'd60856;
        ROM1[69]<=26'd11938; ROM2[69]<=26'd11348; ROM3[69]<=26'd15726; ROM4[69]<=26'd35734;
        ROM1[70]<=26'd19373; ROM2[70]<=26'd18925; ROM3[70]<=26'd30535; ROM4[70]<=26'd64923;
        ROM1[71]<=26'd15362; ROM2[71]<=26'd14975; ROM3[71]<=26'd22541; ROM4[71]<=26'd47339;
        ROM1[72]<=26'd19613; ROM2[72]<=26'd19221; ROM3[72]<=26'd31143; ROM4[72]<=26'd63758;
        ROM1[73]<=26'd16611; ROM2[73]<=26'd16163; ROM3[73]<=26'd25291; ROM4[73]<=26'd50528;
        ROM1[74]<=26'd17726; ROM2[74]<=26'd17192; ROM3[74]<=26'd27712; ROM4[74]<=26'd54247;
        ROM1[75]<=26'd11993; ROM2[75]<=26'd11357; ROM3[75]<=26'd16449; ROM4[75]<=26'd29910;
        ROM1[76]<=26'd13993; ROM2[76]<=26'd13259; ROM3[76]<=26'd20651; ROM4[76]<=26'd37276;
        ROM1[77]<=26'd12685; ROM2[77]<=26'd11874; ROM3[77]<=26'd18212; ROM4[77]<=26'd31037;
        ROM1[78]<=26'd14186; ROM2[78]<=26'd13337; ROM3[78]<=26'd21349; ROM4[78]<=26'd36240;
        ROM1[79]<=26'd12843; ROM2[79]<=26'd12012; ROM3[79]<=26'd18737; ROM4[79]<=26'd29676;
        ROM1[80]<=-26'd1734; ROM2[80]<=-26'd18858; ROM3[80]<=26'd5964; ROM4[80]<=26'd16233;
        ROM1[81]<=-26'd690; ROM2[81]<=-26'd17638; ROM3[81]<=26'd7952; ROM4[81]<=26'd19150;
        ROM1[82]<=-26'd3212; ROM2[82]<=-26'd19883; ROM3[82]<=26'd2698; ROM4[82]<=26'd7257;
        ROM1[83]<=26'd2383; ROM2[83]<=-26'd13898; ROM3[83]<=26'd13558; ROM4[83]<=26'd28431;
        ROM1[84]<=-26'd14473; ROM2[84]<=-26'd22049; ROM3[84]<=-26'd12426; ROM4[84]<=-26'd24655;
        ROM1[85]<=-26'd16262; ROM2[85]<=-26'd23195; ROM3[85]<=-26'd16612; ROM4[85]<=-26'd34241;
        ROM1[86]<=-26'd13346; ROM2[86]<=-26'd19500; ROM3[86]<=-26'd11539; ROM4[86]<=-26'd24799;
        ROM1[87]<=-26'd15932; ROM2[87]<=-26'd21164; ROM3[87]<=-26'd17621; ROM4[87]<=-26'd38182;
        ROM1[88]<=-26'd10922; ROM2[88]<=-26'd15091; ROM3[88]<=-26'd8669; ROM4[88]<=-26'd20696;
        ROM1[89]<=-26'd6837; ROM2[89]<=-26'd9800; ROM3[89]<=-26'd1721; ROM4[89]<=-26'd7273;
        ROM1[90]<=-26'd10523; ROM2[90]<=-26'd12140; ROM3[90]<=-26'd10467; ROM4[90]<=-26'd25977;
        ROM1[91]<=-26'd6226; ROM2[91]<=-26'd6363; ROM3[91]<=-26'd3393; ROM4[91]<=-26'd12208;
        ROM1[92]<=-26'd9059; ROM2[92]<=-26'd7588; ROM3[92]<=-26'd10718; ROM4[92]<=-26'd27913;
        ROM1[93]<=-26'd2608; ROM2[93]<=26'd589; ROM3[93]<=26'd395; ROM4[93]<=-26'd5780;
        ROM1[94]<=-26'd4345; ROM2[94]<=26'd685; ROM3[94]<=-26'd4985; ROM4[94]<=-26'd17424;
        ROM1[95]<=-26'd3368; ROM2[95]<=26'd3589; ROM3[95]<=-26'd5042; ROM4[95]<=-26'd18125;
        ROM1[96]<=-26'd14529; ROM2[96]<=-26'd21947; ROM3[96]<=-26'd13076; ROM4[96]<=-26'd21226;
        ROM1[97]<=-26'd17191; ROM2[97]<=-26'd22536; ROM3[97]<=-26'd20566; ROM4[97]<=-26'd37119;
        ROM1[98]<=-26'd8542; ROM2[98]<=-26'd11766; ROM3[98]<=-26'd5490; ROM4[98]<=-26'd6733;
        ROM1[99]<=-26'd13244; ROM2[99]<=-26'd14315; ROM3[99]<=-26'd17148; ROM4[99]<=-26'd31141;
        ROM1[100]<=26'd10718; ROM2[100]<=26'd3621; ROM3[100]<=26'd20314; ROM4[100]<=26'd43919;
        ROM1[101]<=26'd9436; ROM2[101]<=26'd4500; ROM3[101]<=26'd15486; ROM4[101]<=26'd33514;
        ROM1[102]<=26'd15285; ROM2[102]<=26'd12488; ROM3[102]<=26'd24944; ROM4[102]<=26'd52390;
        ROM1[103]<=26'd19146; ROM2[103]<=26'd18449; ROM3[103]<=26'd30471; ROM4[103]<=26'd63192;
        ROM1[104]<=26'd15252; ROM2[104]<=26'd16596; ROM3[104]<=26'd20549; ROM4[104]<=26'd42304;
        ROM1[105]<=26'd19818; ROM2[105]<=26'd23132; ROM3[105]<=26'd27627; ROM4[105]<=26'd56243;
        ROM1[106]<=26'd21752; ROM2[106]<=26'd26947; ROM3[106]<=26'd29537; ROM4[106]<=26'd59559;
        ROM1[107]<=26'd23302; ROM2[107]<=26'd30277; ROM3[107]<=26'd30788; ROM4[107]<=26'd61493;
        ROM1[108]<=26'd22051; ROM2[108]<=26'd30693; ROM3[108]<=26'd26561; ROM4[108]<=26'd52158;
        ROM1[109]<=26'd29525; ROM2[109]<=26'd39711; ROM3[109]<=26'd39920; ROM4[109]<=26'd78834;
        ROM1[110]<=26'd26761; ROM2[110]<=26'd38359; ROM3[110]<=26'd32945; ROM4[110]<=26'd63782;
        ROM1[111]<=26'd31285; ROM2[111]<=26'd44158; ROM3[111]<=26'd40696; ROM4[111]<=26'd78873;
        ROM1[112]<=26'd14822; ROM2[112]<=26'd12445; ROM3[112]<=26'd23011; ROM4[112]<=26'd55701;
        ROM1[113]<=26'd12524; ROM2[113]<=26'd11138; ROM3[113]<=26'd17426; ROM4[113]<=26'd43362;
        ROM1[114]<=26'd17619; ROM2[114]<=26'd17082; ROM3[114]<=26'd26785; ROM4[114]<=26'd61610;
        ROM1[115]<=26'd14940; ROM2[115]<=26'd15113; ROM3[115]<=26'd20746; ROM4[115]<=26'd48247;
        ROM1[116]<=26'd19527; ROM2[116]<=26'd20275; ROM3[116]<=26'd29385; ROM4[116]<=26'd64932;
        ROM1[117]<=26'd1188; ROM2[117]<=26'd10578; ROM3[117]<=26'd505; ROM4[117]<=26'd5888;
        ROM1[118]<=26'd4045; ROM2[118]<=26'd13765; ROM3[118]<=26'd5950; ROM4[118]<=26'd15943;
        ROM1[119]<=26'd2793; ROM2[119]<=26'd12738; ROM3[119]<=26'd3295; ROM4[119]<=26'd9359;
        ROM1[120]<=26'd3274; ROM2[120]<=26'd13349; ROM3[120]<=26'd4207; ROM4[120]<=26'd10058;
        ROM1[121]<=26'd1580; ROM2[121]<=26'd11707; ROM3[121]<=26'd857; ROM4[121]<=26'd1992;
        ROM1[122]<=26'd5388; ROM2[122]<=26'd15502; ROM3[122]<=26'd8581; ROM4[122]<=26'd16605;
        ROM1[123]<=26'd2870; ROM2[123]<=26'd12925; ROM3[123]<=26'd3705; ROM4[123]<=26'd5376;
        ROM1[124]<=26'd1079; ROM2[124]<=26'd11044; ROM3[124]<=26'd315; ROM4[124]<=-26'd2819;
        ROM1[125]<=26'd2575; ROM2[125]<=26'd12438; ROM3[125]<=26'd3513; ROM4[125]<=26'd2488;
        ROM1[126]<=-26'd2229; ROM2[126]<=26'd7538; ROM3[126]<=-26'd5897; ROM4[126]<=-26'd18048;
        ROM1[127]<=-26'd16272; ROM2[127]<=-26'd22962; ROM3[127]<=-26'd17426; ROM4[127]<=-26'd28994;
	end
	else begin
		if(cnt == 7'd127) begin
				cnt<=0;
			end
		//?��?��?�� addr?��?��.
		data1 <= ROM1[cnt];
		data2 <= ROM2[cnt];
		data3 <= ROM3[cnt];
		data4 <= ROM4[cnt];
		cnt <= cnt+1'b1;
	end
end
endmodule 
