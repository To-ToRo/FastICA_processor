//출처 : https://verilogguide.readthedocs.io/en/latest/verilog/designs.html#read-only-memory-rom

module ROM(
    input wire clk,
	input wire En,
    input wire  [13:0] addr,
    output reg unsigned [25:0] data1,
	output reg unsigned [25:0] data2,
	output reg unsigned [25:0] data3,
	output reg unsigned [25:0] data4
);

//ROM[0]의 크기 : 16bit(한 시그널의 크기) * 4(4개의 시그널) 
// 각각의 시그널이 총 1000sample이 있으므로 addr은  16비트로 표현(0~39999 < 0~65536) 

reg unsigned [25:0] ROM1[0:9999];
reg unsigned [25:0] ROM2[0:9999];
reg unsigned [25:0] ROM3[0:9999];
reg unsigned [25:0] ROM4[0:9999];
reg [6:0] cnt;

always @(posedge clk) begin
	if(!En) begin
		cnt<=0;
data1<=0;
data2<=0;
data3<=0;
data4<=0;

ROM1[0]<=26'd1961154; ROM2[0]<=26'd11295750; ROM3[0]<=26'd9760920; ROM4[0]<=26'd23462602;
ROM1[1]<=26'd1962156; ROM2[1]<=26'd11296488; ROM3[1]<=26'd9764935; ROM4[1]<=26'd23465762;
ROM1[2]<=26'd1951852; ROM2[2]<=26'd11292489; ROM3[2]<=26'd9764653; ROM4[2]<=26'd23464634;
ROM1[3]<=26'd1937555; ROM2[3]<=26'd11282542; ROM3[3]<=26'd9758485; ROM4[3]<=26'd23455973;
ROM1[4]<=26'd1932118; ROM2[4]<=26'd11279931; ROM3[4]<=26'd9758040; ROM4[4]<=26'd23455320;
ROM1[5]<=26'd1927580; ROM2[5]<=26'd11279516; ROM3[5]<=26'd9759644; ROM4[5]<=26'd23454723;
ROM1[6]<=26'd1932145; ROM2[6]<=26'd11284885; ROM3[6]<=26'd9763797; ROM4[6]<=26'd23458732;
ROM1[7]<=26'd1938850; ROM2[7]<=26'd11285707; ROM3[7]<=26'd9757271; ROM4[7]<=26'd23456575;
ROM1[8]<=26'd1942834; ROM2[8]<=26'd11278973; ROM3[8]<=26'd9743882; ROM4[8]<=26'd23448230;
ROM1[9]<=26'd1947999; ROM2[9]<=26'd11280626; ROM3[9]<=26'd9743229; ROM4[9]<=26'd23449963;
ROM1[10]<=26'd1943279; ROM2[10]<=26'd11280461; ROM3[10]<=26'd9745995; ROM4[10]<=26'd23451243;
ROM1[11]<=26'd1939937; ROM2[11]<=26'd11281789; ROM3[11]<=26'd9753958; ROM4[11]<=26'd23455867;
ROM1[12]<=26'd1935994; ROM2[12]<=26'd11282627; ROM3[12]<=26'd9757700; ROM4[12]<=26'd23458109;
ROM1[13]<=26'd1924973; ROM2[13]<=26'd11277722; ROM3[13]<=26'd9755802; ROM4[13]<=26'd23454760;
ROM1[14]<=26'd1919812; ROM2[14]<=26'd11274650; ROM3[14]<=26'd9753633; ROM4[14]<=26'd23450160;
ROM1[15]<=26'd1927410; ROM2[15]<=26'd11278690; ROM3[15]<=26'd9751149; ROM4[15]<=26'd23450337;
ROM1[16]<=26'd1947915; ROM2[16]<=26'd11289330; ROM3[16]<=26'd9754069; ROM4[16]<=26'd23457957;
ROM1[17]<=26'd1959909; ROM2[17]<=26'd11293804; ROM3[17]<=26'd9754082; ROM4[17]<=26'd23462277;
ROM1[18]<=26'd1950663; ROM2[18]<=26'd11285517; ROM3[18]<=26'd9745105; ROM4[18]<=26'd23454720;
ROM1[19]<=26'd1937432; ROM2[19]<=26'd11281118; ROM3[19]<=26'd9743059; ROM4[19]<=26'd23449931;
ROM1[20]<=26'd1930425; ROM2[20]<=26'd11279268; ROM3[20]<=26'd9745252; ROM4[20]<=26'd23446984;
ROM1[21]<=26'd1923426; ROM2[21]<=26'd11275870; ROM3[21]<=26'd9742941; ROM4[21]<=26'd23441554;
ROM1[22]<=26'd1919051; ROM2[22]<=26'd11277509; ROM3[22]<=26'd9744980; ROM4[22]<=26'd23444016;
ROM1[23]<=26'd1922878; ROM2[23]<=26'd11280124; ROM3[23]<=26'd9744453; ROM4[23]<=26'd23445806;
ROM1[24]<=26'd1932339; ROM2[24]<=26'd11280163; ROM3[24]<=26'd9737673; ROM4[24]<=26'd23442634;
ROM1[25]<=26'd1943529; ROM2[25]<=26'd11281605; ROM3[25]<=26'd9731070; ROM4[25]<=26'd23442249;
ROM1[26]<=26'd1944965; ROM2[26]<=26'd11283599; ROM3[26]<=26'd9731145; ROM4[26]<=26'd23443506;
ROM1[27]<=26'd1938494; ROM2[27]<=26'd11282705; ROM3[27]<=26'd9733700; ROM4[27]<=26'd23443026;
ROM1[28]<=26'd1929589; ROM2[28]<=26'd11282125; ROM3[28]<=26'd9737100; ROM4[28]<=26'd23442595;
ROM1[29]<=26'd1921593; ROM2[29]<=26'd11280934; ROM3[29]<=26'd9737668; ROM4[29]<=26'd23441334;
ROM1[30]<=26'd1916748; ROM2[30]<=26'd11281545; ROM3[30]<=26'd9737858; ROM4[30]<=26'd23441265;
ROM1[31]<=26'd1921909; ROM2[31]<=26'd11284469; ROM3[31]<=26'd9739903; ROM4[31]<=26'd23443256;
ROM1[32]<=26'd1934859; ROM2[32]<=26'd11288100; ROM3[32]<=26'd9739189; ROM4[32]<=26'd23447065;
ROM1[33]<=26'd1949417; ROM2[33]<=26'd11291144; ROM3[33]<=26'd9736336; ROM4[33]<=26'd23450499;
ROM1[34]<=26'd1951585; ROM2[34]<=26'd11290860; ROM3[34]<=26'd9738574; ROM4[34]<=26'd23452905;
ROM1[35]<=26'd1945722; ROM2[35]<=26'd11291359; ROM3[35]<=26'd9743956; ROM4[35]<=26'd23455870;
ROM1[36]<=26'd1941165; ROM2[36]<=26'd11293078; ROM3[36]<=26'd9750541; ROM4[36]<=26'd23458048;
ROM1[37]<=26'd1939567; ROM2[37]<=26'd11296686; ROM3[37]<=26'd9756049; ROM4[37]<=26'd23457640;
ROM1[38]<=26'd1938652; ROM2[38]<=26'd11301078; ROM3[38]<=26'd9759598; ROM4[38]<=26'd23458656;
ROM1[39]<=26'd1936479; ROM2[39]<=26'd11298737; ROM3[39]<=26'd9759258; ROM4[39]<=26'd23456974;
ROM1[40]<=26'd1943079; ROM2[40]<=26'd11298651; ROM3[40]<=26'd9758649; ROM4[40]<=26'd23458328;
ROM1[41]<=26'd1949436; ROM2[41]<=26'd11292299; ROM3[41]<=26'd9748022; ROM4[41]<=26'd23452512;
ROM1[42]<=26'd1950769; ROM2[42]<=26'd11285642; ROM3[42]<=26'd9738145; ROM4[42]<=26'd23446462;
ROM1[43]<=26'd1948502; ROM2[43]<=26'd11285707; ROM3[43]<=26'd9739814; ROM4[43]<=26'd23446068;
ROM1[44]<=26'd1941389; ROM2[44]<=26'd11285027; ROM3[44]<=26'd9742663; ROM4[44]<=26'd23445456;
ROM1[45]<=26'd1933402; ROM2[45]<=26'd11284643; ROM3[45]<=26'd9745262; ROM4[45]<=26'd23447312;
ROM1[46]<=26'd1928631; ROM2[46]<=26'd11283994; ROM3[46]<=26'd9746762; ROM4[46]<=26'd23446792;
ROM1[47]<=26'd1925463; ROM2[47]<=26'd11285381; ROM3[47]<=26'd9746387; ROM4[47]<=26'd23445621;
ROM1[48]<=26'd1929631; ROM2[48]<=26'd11286935; ROM3[48]<=26'd9747127; ROM4[48]<=26'd23448121;
ROM1[49]<=26'd1940649; ROM2[49]<=26'd11288846; ROM3[49]<=26'd9744545; ROM4[49]<=26'd23448989;
ROM1[50]<=26'd1948831; ROM2[50]<=26'd11289571; ROM3[50]<=26'd9739535; ROM4[50]<=26'd23446325;
ROM1[51]<=26'd1952167; ROM2[51]<=26'd11295557; ROM3[51]<=26'd9744038; ROM4[51]<=26'd23452021;
ROM1[52]<=26'd1942909; ROM2[52]<=26'd11294197; ROM3[52]<=26'd9742828; ROM4[52]<=26'd23451432;
ROM1[53]<=26'd1930296; ROM2[53]<=26'd11285206; ROM3[53]<=26'd9738079; ROM4[53]<=26'd23442719;
ROM1[54]<=26'd1929219; ROM2[54]<=26'd11286382; ROM3[54]<=26'd9743426; ROM4[54]<=26'd23445080;
ROM1[55]<=26'd1925317; ROM2[55]<=26'd11287228; ROM3[55]<=26'd9747592; ROM4[55]<=26'd23446912;
ROM1[56]<=26'd1923085; ROM2[56]<=26'd11284804; ROM3[56]<=26'd9745116; ROM4[56]<=26'd23443392;
ROM1[57]<=26'd1934691; ROM2[57]<=26'd11289600; ROM3[57]<=26'd9744981; ROM4[57]<=26'd23445443;
ROM1[58]<=26'd1949080; ROM2[58]<=26'd11292049; ROM3[58]<=26'd9740619; ROM4[58]<=26'd23446350;
ROM1[59]<=26'd1950525; ROM2[59]<=26'd11289127; ROM3[59]<=26'd9736845; ROM4[59]<=26'd23445848;
ROM1[60]<=26'd1945336; ROM2[60]<=26'd11289807; ROM3[60]<=26'd9740891; ROM4[60]<=26'd23447309;
ROM1[61]<=26'd1944937; ROM2[61]<=26'd11294842; ROM3[61]<=26'd9753120; ROM4[61]<=26'd23456142;
ROM1[62]<=26'd1946431; ROM2[62]<=26'd11300540; ROM3[62]<=26'd9764014; ROM4[62]<=26'd23465083;
ROM1[63]<=26'd1936483; ROM2[63]<=26'd11294196; ROM3[63]<=26'd9762270; ROM4[63]<=26'd23459563;
ROM1[64]<=26'd1930949; ROM2[64]<=26'd11289243; ROM3[64]<=26'd9758967; ROM4[64]<=26'd23455561;
ROM1[65]<=26'd1936621; ROM2[65]<=26'd11288950; ROM3[65]<=26'd9757594; ROM4[65]<=26'd23455858;
ROM1[66]<=26'd1946582; ROM2[66]<=26'd11285961; ROM3[66]<=26'd9750838; ROM4[66]<=26'd23454158;
ROM1[67]<=26'd1954454; ROM2[67]<=26'd11286942; ROM3[67]<=26'd9748385; ROM4[67]<=26'd23456209;
ROM1[68]<=26'd1953657; ROM2[68]<=26'd11287241; ROM3[68]<=26'd9751178; ROM4[68]<=26'd23457816;
ROM1[69]<=26'd1946212; ROM2[69]<=26'd11285860; ROM3[69]<=26'd9754499; ROM4[69]<=26'd23457459;
ROM1[70]<=26'd1939077; ROM2[70]<=26'd11285181; ROM3[70]<=26'd9758223; ROM4[70]<=26'd23457458;
ROM1[71]<=26'd1938722; ROM2[71]<=26'd11288200; ROM3[71]<=26'd9764886; ROM4[71]<=26'd23461460;
ROM1[72]<=26'd1937317; ROM2[72]<=26'd11290100; ROM3[72]<=26'd9767954; ROM4[72]<=26'd23463635;
ROM1[73]<=26'd1939191; ROM2[73]<=26'd11290674; ROM3[73]<=26'd9763869; ROM4[73]<=26'd23462185;
ROM1[74]<=26'd1944954; ROM2[74]<=26'd11288617; ROM3[74]<=26'd9753847; ROM4[74]<=26'd23457195;
ROM1[75]<=26'd1949629; ROM2[75]<=26'd11284668; ROM3[75]<=26'd9741066; ROM4[75]<=26'd23449224;
ROM1[76]<=26'd1945987; ROM2[76]<=26'd11281152; ROM3[76]<=26'd9735773; ROM4[76]<=26'd23444384;
ROM1[77]<=26'd1941151; ROM2[77]<=26'd11282905; ROM3[77]<=26'd9740152; ROM4[77]<=26'd23447438;
ROM1[78]<=26'd1939326; ROM2[78]<=26'd11287744; ROM3[78]<=26'd9749697; ROM4[78]<=26'd23454555;
ROM1[79]<=26'd1929841; ROM2[79]<=26'd11284647; ROM3[79]<=26'd9748884; ROM4[79]<=26'd23450622;
ROM1[80]<=26'd1922903; ROM2[80]<=26'd11281496; ROM3[80]<=26'd9747492; ROM4[80]<=26'd23448932;
ROM1[81]<=26'd1921634; ROM2[81]<=26'd11279095; ROM3[81]<=26'd9744887; ROM4[81]<=26'd23447496;
ROM1[82]<=26'd1925923; ROM2[82]<=26'd11276516; ROM3[82]<=26'd9734485; ROM4[82]<=26'd23439240;
ROM1[83]<=26'd1938662; ROM2[83]<=26'd11278855; ROM3[83]<=26'd9728967; ROM4[83]<=26'd23438824;
ROM1[84]<=26'd1943159; ROM2[84]<=26'd11281594; ROM3[84]<=26'd9730029; ROM4[84]<=26'd23442357;
ROM1[85]<=26'd1939924; ROM2[85]<=26'd11285152; ROM3[85]<=26'd9734082; ROM4[85]<=26'd23444438;
ROM1[86]<=26'd1932039; ROM2[86]<=26'd11284987; ROM3[86]<=26'd9735880; ROM4[86]<=26'd23442662;
ROM1[87]<=26'd1929620; ROM2[87]<=26'd11286757; ROM3[87]<=26'd9739044; ROM4[87]<=26'd23444328;
ROM1[88]<=26'd1924225; ROM2[88]<=26'd11288743; ROM3[88]<=26'd9743039; ROM4[88]<=26'd23445026;
ROM1[89]<=26'd1916973; ROM2[89]<=26'd11283282; ROM3[89]<=26'd9738115; ROM4[89]<=26'd23437990;
ROM1[90]<=26'd1922575; ROM2[90]<=26'd11283540; ROM3[90]<=26'd9737387; ROM4[90]<=26'd23439251;
ROM1[91]<=26'd1936296; ROM2[91]<=26'd11286817; ROM3[91]<=26'd9734723; ROM4[91]<=26'd23442685;
ROM1[92]<=26'd1939584; ROM2[92]<=26'd11283422; ROM3[92]<=26'd9726503; ROM4[92]<=26'd23436941;
ROM1[93]<=26'd1937164; ROM2[93]<=26'd11283500; ROM3[93]<=26'd9726965; ROM4[93]<=26'd23437455;
ROM1[94]<=26'd1932322; ROM2[94]<=26'd11285781; ROM3[94]<=26'd9733560; ROM4[94]<=26'd23441496;
ROM1[95]<=26'd1920488; ROM2[95]<=26'd11278700; ROM3[95]<=26'd9731846; ROM4[95]<=26'd23436698;
ROM1[96]<=26'd1916942; ROM2[96]<=26'd11280434; ROM3[96]<=26'd9736033; ROM4[96]<=26'd23439187;
ROM1[97]<=26'd1920533; ROM2[97]<=26'd11288262; ROM3[97]<=26'd9746560; ROM4[97]<=26'd23446882;
ROM1[98]<=26'd1925831; ROM2[98]<=26'd11288867; ROM3[98]<=26'd9746445; ROM4[98]<=26'd23448734;
ROM1[99]<=26'd1931810; ROM2[99]<=26'd11286281; ROM3[99]<=26'd9739158; ROM4[99]<=26'd23445175;
ROM1[100]<=26'd1937615; ROM2[100]<=26'd11283678; ROM3[100]<=26'd9729007; ROM4[100]<=26'd23439241;
ROM1[101]<=26'd1933919; ROM2[101]<=26'd11279713; ROM3[101]<=26'd9724752; ROM4[101]<=26'd23436104;
ROM1[102]<=26'd1923364; ROM2[102]<=26'd11275261; ROM3[102]<=26'd9722862; ROM4[102]<=26'd23432566;
ROM1[103]<=26'd1921435; ROM2[103]<=26'd11277817; ROM3[103]<=26'd9729910; ROM4[103]<=26'd23434950;
ROM1[104]<=26'd1921794; ROM2[104]<=26'd11278409; ROM3[104]<=26'd9734989; ROM4[104]<=26'd23439083;
ROM1[105]<=26'd1915409; ROM2[105]<=26'd11275035; ROM3[105]<=26'd9734000; ROM4[105]<=26'd23436421;
ROM1[106]<=26'd1917585; ROM2[106]<=26'd11276014; ROM3[106]<=26'd9733833; ROM4[106]<=26'd23435452;
ROM1[107]<=26'd1931223; ROM2[107]<=26'd11281967; ROM3[107]<=26'd9735592; ROM4[107]<=26'd23441917;
ROM1[108]<=26'd1946777; ROM2[108]<=26'd11288424; ROM3[108]<=26'd9736396; ROM4[108]<=26'd23446919;
ROM1[109]<=26'd1948677; ROM2[109]<=26'd11289711; ROM3[109]<=26'd9734753; ROM4[109]<=26'd23447325;
ROM1[110]<=26'd1943760; ROM2[110]<=26'd11288559; ROM3[110]<=26'd9737535; ROM4[110]<=26'd23448833;
ROM1[111]<=26'd1938847; ROM2[111]<=26'd11287408; ROM3[111]<=26'd9742876; ROM4[111]<=26'd23449971;
ROM1[112]<=26'd1937798; ROM2[112]<=26'd11289693; ROM3[112]<=26'd9750810; ROM4[112]<=26'd23454260;
ROM1[113]<=26'd1932864; ROM2[113]<=26'd11290497; ROM3[113]<=26'd9753981; ROM4[113]<=26'd23455126;
ROM1[114]<=26'd1925784; ROM2[114]<=26'd11285357; ROM3[114]<=26'd9749152; ROM4[114]<=26'd23450241;
ROM1[115]<=26'd1929057; ROM2[115]<=26'd11283819; ROM3[115]<=26'd9745611; ROM4[115]<=26'd23447666;
ROM1[116]<=26'd1942090; ROM2[116]<=26'd11283575; ROM3[116]<=26'd9740930; ROM4[116]<=26'd23445625;
ROM1[117]<=26'd1954432; ROM2[117]<=26'd11283857; ROM3[117]<=26'd9740276; ROM4[117]<=26'd23447606;
ROM1[118]<=26'd1957779; ROM2[118]<=26'd11289375; ROM3[118]<=26'd9747203; ROM4[118]<=26'd23453797;
ROM1[119]<=26'd1950954; ROM2[119]<=26'd11289068; ROM3[119]<=26'd9751227; ROM4[119]<=26'd23456637;
ROM1[120]<=26'd1943095; ROM2[120]<=26'd11288813; ROM3[120]<=26'd9753092; ROM4[120]<=26'd23458179;
ROM1[121]<=26'd1939229; ROM2[121]<=26'd11290848; ROM3[121]<=26'd9758201; ROM4[121]<=26'd23461077;
ROM1[122]<=26'd1944604; ROM2[122]<=26'd11297460; ROM3[122]<=26'd9768077; ROM4[122]<=26'd23469461;
ROM1[123]<=26'd1949157; ROM2[123]<=26'd11298374; ROM3[123]<=26'd9763990; ROM4[123]<=26'd23469280;
ROM1[124]<=26'd1951370; ROM2[124]<=26'd11287473; ROM3[124]<=26'd9748087; ROM4[124]<=26'd23457432;
ROM1[125]<=26'd1955665; ROM2[125]<=26'd11279086; ROM3[125]<=26'd9735977; ROM4[125]<=26'd23451406;
ROM1[126]<=26'd1949627; ROM2[126]<=26'd11274542; ROM3[126]<=26'd9731743; ROM4[126]<=26'd23448339;
ROM1[127]<=26'd1946214; ROM2[127]<=26'd11277978; ROM3[127]<=26'd9738813; ROM4[127]<=26'd23450520;
ROM1[128]<=26'd1940502; ROM2[128]<=26'd11278635; ROM3[128]<=26'd9744835; ROM4[128]<=26'd23453446;
ROM1[129]<=26'd1933802; ROM2[129]<=26'd11276416; ROM3[129]<=26'd9746462; ROM4[129]<=26'd23451895;
ROM1[130]<=26'd1926431; ROM2[130]<=26'd11273631; ROM3[130]<=26'd9746270; ROM4[130]<=26'd23448534;
ROM1[131]<=26'd1925104; ROM2[131]<=26'd11270381; ROM3[131]<=26'd9746259; ROM4[131]<=26'd23447309;
ROM1[132]<=26'd1934760; ROM2[132]<=26'd11273884; ROM3[132]<=26'd9746602; ROM4[132]<=26'd23448833;
ROM1[133]<=26'd1947158; ROM2[133]<=26'd11279211; ROM3[133]<=26'd9744271; ROM4[133]<=26'd23451517;
ROM1[134]<=26'd1951226; ROM2[134]<=26'd11282453; ROM3[134]<=26'd9744106; ROM4[134]<=26'd23452896;
ROM1[135]<=26'd1944462; ROM2[135]<=26'd11281949; ROM3[135]<=26'd9746136; ROM4[135]<=26'd23452207;
ROM1[136]<=26'd1932940; ROM2[136]<=26'd11276417; ROM3[136]<=26'd9745569; ROM4[136]<=26'd23447872;
ROM1[137]<=26'd1924728; ROM2[137]<=26'd11272973; ROM3[137]<=26'd9744558; ROM4[137]<=26'd23442850;
ROM1[138]<=26'd1911343; ROM2[138]<=26'd11267613; ROM3[138]<=26'd9742053; ROM4[138]<=26'd23438120;
ROM1[139]<=26'd1907384; ROM2[139]<=26'd11267595; ROM3[139]<=26'd9740517; ROM4[139]<=26'd23436997;
ROM1[140]<=26'd1920364; ROM2[140]<=26'd11277231; ROM3[140]<=26'd9744060; ROM4[140]<=26'd23444418;
ROM1[141]<=26'd1945318; ROM2[141]<=26'd11290980; ROM3[141]<=26'd9750702; ROM4[141]<=26'd23457347;
ROM1[142]<=26'd1956568; ROM2[142]<=26'd11295029; ROM3[142]<=26'd9751079; ROM4[142]<=26'd23462133;
ROM1[143]<=26'd1946378; ROM2[143]<=26'd11288668; ROM3[143]<=26'd9744715; ROM4[143]<=26'd23455062;
ROM1[144]<=26'd1935464; ROM2[144]<=26'd11284761; ROM3[144]<=26'd9742824; ROM4[144]<=26'd23451410;
ROM1[145]<=26'd1919186; ROM2[145]<=26'd11273033; ROM3[145]<=26'd9736302; ROM4[145]<=26'd23440604;
ROM1[146]<=26'd1908112; ROM2[146]<=26'd11264226; ROM3[146]<=26'd9732258; ROM4[146]<=26'd23433134;
ROM1[147]<=26'd1906386; ROM2[147]<=26'd11264751; ROM3[147]<=26'd9734290; ROM4[147]<=26'd23434762;
ROM1[148]<=26'd1908286; ROM2[148]<=26'd11266231; ROM3[148]<=26'd9732885; ROM4[148]<=26'd23435141;
ROM1[149]<=26'd1918318; ROM2[149]<=26'd11267789; ROM3[149]<=26'd9726921; ROM4[149]<=26'd23434255;
ROM1[150]<=26'd1927631; ROM2[150]<=26'd11267369; ROM3[150]<=26'd9719561; ROM4[150]<=26'd23429853;
ROM1[151]<=26'd1927947; ROM2[151]<=26'd11268565; ROM3[151]<=26'd9722544; ROM4[151]<=26'd23431628;
ROM1[152]<=26'd1921895; ROM2[152]<=26'd11268372; ROM3[152]<=26'd9727969; ROM4[152]<=26'd23432688;
ROM1[153]<=26'd1911211; ROM2[153]<=26'd11265171; ROM3[153]<=26'd9729701; ROM4[153]<=26'd23430445;
ROM1[154]<=26'd1908001; ROM2[154]<=26'd11268053; ROM3[154]<=26'd9734679; ROM4[154]<=26'd23434732;
ROM1[155]<=26'd1907994; ROM2[155]<=26'd11271745; ROM3[155]<=26'd9741482; ROM4[155]<=26'd23437710;
ROM1[156]<=26'd1913404; ROM2[156]<=26'd11275940; ROM3[156]<=26'd9743814; ROM4[156]<=26'd23440062;
ROM1[157]<=26'd1928777; ROM2[157]<=26'd11284237; ROM3[157]<=26'd9745744; ROM4[157]<=26'd23445390;
ROM1[158]<=26'd1941889; ROM2[158]<=26'd11283626; ROM3[158]<=26'd9740097; ROM4[158]<=26'd23442837;
ROM1[159]<=26'd1942239; ROM2[159]<=26'd11280407; ROM3[159]<=26'd9734513; ROM4[159]<=26'd23440094;
ROM1[160]<=26'd1936134; ROM2[160]<=26'd11280166; ROM3[160]<=26'd9735252; ROM4[160]<=26'd23439961;
ROM1[161]<=26'd1927847; ROM2[161]<=26'd11278836; ROM3[161]<=26'd9737104; ROM4[161]<=26'd23439491;
ROM1[162]<=26'd1922779; ROM2[162]<=26'd11278055; ROM3[162]<=26'd9738264; ROM4[162]<=26'd23440134;
ROM1[163]<=26'd1920461; ROM2[163]<=26'd11280884; ROM3[163]<=26'd9743930; ROM4[163]<=26'd23442346;
ROM1[164]<=26'd1921354; ROM2[164]<=26'd11282948; ROM3[164]<=26'd9746466; ROM4[164]<=26'd23444309;
ROM1[165]<=26'd1929882; ROM2[165]<=26'd11285370; ROM3[165]<=26'd9744475; ROM4[165]<=26'd23444854;
ROM1[166]<=26'd1942822; ROM2[166]<=26'd11288367; ROM3[166]<=26'd9742400; ROM4[166]<=26'd23444880;
ROM1[167]<=26'd1947750; ROM2[167]<=26'd11287549; ROM3[167]<=26'd9735562; ROM4[167]<=26'd23442331;
ROM1[168]<=26'd1946762; ROM2[168]<=26'd11290237; ROM3[168]<=26'd9738855; ROM4[168]<=26'd23444941;
ROM1[169]<=26'd1941569; ROM2[169]<=26'd11290595; ROM3[169]<=26'd9742980; ROM4[169]<=26'd23445592;
ROM1[170]<=26'd1930025; ROM2[170]<=26'd11286186; ROM3[170]<=26'd9738858; ROM4[170]<=26'd23439575;
ROM1[171]<=26'd1922408; ROM2[171]<=26'd11281696; ROM3[171]<=26'd9737504; ROM4[171]<=26'd23437648;
ROM1[172]<=26'd1919532; ROM2[172]<=26'd11279357; ROM3[172]<=26'd9738583; ROM4[172]<=26'd23436988;
ROM1[173]<=26'd1928782; ROM2[173]<=26'd11283984; ROM3[173]<=26'd9742828; ROM4[173]<=26'd23443472;
ROM1[174]<=26'd1944382; ROM2[174]<=26'd11286503; ROM3[174]<=26'd9741423; ROM4[174]<=26'd23444839;
ROM1[175]<=26'd1954104; ROM2[175]<=26'd11285833; ROM3[175]<=26'd9735742; ROM4[175]<=26'd23442856;
ROM1[176]<=26'd1950731; ROM2[176]<=26'd11281644; ROM3[176]<=26'd9731711; ROM4[176]<=26'd23441252;
ROM1[177]<=26'd1939840; ROM2[177]<=26'd11277370; ROM3[177]<=26'd9731170; ROM4[177]<=26'd23438600;
ROM1[178]<=26'd1933585; ROM2[178]<=26'd11278721; ROM3[178]<=26'd9736702; ROM4[178]<=26'd23441704;
ROM1[179]<=26'd1929998; ROM2[179]<=26'd11281333; ROM3[179]<=26'd9741653; ROM4[179]<=26'd23445912;
ROM1[180]<=26'd1925166; ROM2[180]<=26'd11281057; ROM3[180]<=26'd9744334; ROM4[180]<=26'd23445427;
ROM1[181]<=26'd1925234; ROM2[181]<=26'd11278828; ROM3[181]<=26'd9741364; ROM4[181]<=26'd23441025;
ROM1[182]<=26'd1937165; ROM2[182]<=26'd11280590; ROM3[182]<=26'd9739633; ROM4[182]<=26'd23444451;
ROM1[183]<=26'd1955009; ROM2[183]<=26'd11286965; ROM3[183]<=26'd9739854; ROM4[183]<=26'd23449224;
ROM1[184]<=26'd1956287; ROM2[184]<=26'd11288155; ROM3[184]<=26'd9737753; ROM4[184]<=26'd23448910;
ROM1[185]<=26'd1943774; ROM2[185]<=26'd11283124; ROM3[185]<=26'd9734273; ROM4[185]<=26'd23446091;
ROM1[186]<=26'd1933153; ROM2[186]<=26'd11280418; ROM3[186]<=26'd9736411; ROM4[186]<=26'd23445112;
ROM1[187]<=26'd1926498; ROM2[187]<=26'd11279752; ROM3[187]<=26'd9738446; ROM4[187]<=26'd23444705;
ROM1[188]<=26'd1927686; ROM2[188]<=26'd11288586; ROM3[188]<=26'd9746929; ROM4[188]<=26'd23450803;
ROM1[189]<=26'd1929452; ROM2[189]<=26'd11293300; ROM3[189]<=26'd9753684; ROM4[189]<=26'd23454037;
ROM1[190]<=26'd1925486; ROM2[190]<=26'd11285896; ROM3[190]<=26'd9744165; ROM4[190]<=26'd23446229;
ROM1[191]<=26'd1934985; ROM2[191]<=26'd11285098; ROM3[191]<=26'd9736717; ROM4[191]<=26'd23443432;
ROM1[192]<=26'd1942388; ROM2[192]<=26'd11283467; ROM3[192]<=26'd9732617; ROM4[192]<=26'd23442576;
ROM1[193]<=26'd1936947; ROM2[193]<=26'd11281030; ROM3[193]<=26'd9730565; ROM4[193]<=26'd23441687;
ROM1[194]<=26'd1936352; ROM2[194]<=26'd11288839; ROM3[194]<=26'd9739565; ROM4[194]<=26'd23447536;
ROM1[195]<=26'd1929882; ROM2[195]<=26'd11287872; ROM3[195]<=26'd9743077; ROM4[195]<=26'd23447666;
ROM1[196]<=26'd1913888; ROM2[196]<=26'd11277812; ROM3[196]<=26'd9737302; ROM4[196]<=26'd23439442;
ROM1[197]<=26'd1909669; ROM2[197]<=26'd11277261; ROM3[197]<=26'd9739398; ROM4[197]<=26'd23438286;
ROM1[198]<=26'd1920359; ROM2[198]<=26'd11282384; ROM3[198]<=26'd9742923; ROM4[198]<=26'd23442910;
ROM1[199]<=26'd1936897; ROM2[199]<=26'd11287463; ROM3[199]<=26'd9742652; ROM4[199]<=26'd23447498;
ROM1[200]<=26'd1945169; ROM2[200]<=26'd11287702; ROM3[200]<=26'd9737254; ROM4[200]<=26'd23447305;
ROM1[201]<=26'd1939192; ROM2[201]<=26'd11281851; ROM3[201]<=26'd9732118; ROM4[201]<=26'd23442269;
ROM1[202]<=26'd1930484; ROM2[202]<=26'd11277748; ROM3[202]<=26'd9731566; ROM4[202]<=26'd23440399;
ROM1[203]<=26'd1921809; ROM2[203]<=26'd11274464; ROM3[203]<=26'd9732890; ROM4[203]<=26'd23438930;
ROM1[204]<=26'd1917912; ROM2[204]<=26'd11274681; ROM3[204]<=26'd9735524; ROM4[204]<=26'd23438808;
ROM1[205]<=26'd1915813; ROM2[205]<=26'd11278573; ROM3[205]<=26'd9740332; ROM4[205]<=26'd23442466;
ROM1[206]<=26'd1916361; ROM2[206]<=26'd11281450; ROM3[206]<=26'd9741246; ROM4[206]<=26'd23443629;
ROM1[207]<=26'd1923565; ROM2[207]<=26'd11281336; ROM3[207]<=26'd9736225; ROM4[207]<=26'd23442637;
ROM1[208]<=26'd1936121; ROM2[208]<=26'd11282183; ROM3[208]<=26'd9732152; ROM4[208]<=26'd23443538;
ROM1[209]<=26'd1939252; ROM2[209]<=26'd11282760; ROM3[209]<=26'd9730643; ROM4[209]<=26'd23442760;
ROM1[210]<=26'd1934413; ROM2[210]<=26'd11280983; ROM3[210]<=26'd9732080; ROM4[210]<=26'd23442571;
ROM1[211]<=26'd1926752; ROM2[211]<=26'd11279076; ROM3[211]<=26'd9734428; ROM4[211]<=26'd23441520;
ROM1[212]<=26'd1922796; ROM2[212]<=26'd11278565; ROM3[212]<=26'd9734860; ROM4[212]<=26'd23441283;
ROM1[213]<=26'd1917512; ROM2[213]<=26'd11277411; ROM3[213]<=26'd9738552; ROM4[213]<=26'd23443125;
ROM1[214]<=26'd1913388; ROM2[214]<=26'd11276163; ROM3[214]<=26'd9738591; ROM4[214]<=26'd23443512;
ROM1[215]<=26'd1919009; ROM2[215]<=26'd11276606; ROM3[215]<=26'd9734473; ROM4[215]<=26'd23442090;
ROM1[216]<=26'd1937566; ROM2[216]<=26'd11282568; ROM3[216]<=26'd9732267; ROM4[216]<=26'd23443669;
ROM1[217]<=26'd1953891; ROM2[217]<=26'd11292928; ROM3[217]<=26'd9735129; ROM4[217]<=26'd23452410;
ROM1[218]<=26'd1949110; ROM2[218]<=26'd11291650; ROM3[218]<=26'd9735356; ROM4[218]<=26'd23451970;
ROM1[219]<=26'd1939398; ROM2[219]<=26'd11288416; ROM3[219]<=26'd9737243; ROM4[219]<=26'd23449437;
ROM1[220]<=26'd1931090; ROM2[220]<=26'd11284245; ROM3[220]<=26'd9738734; ROM4[220]<=26'd23448479;
ROM1[221]<=26'd1919647; ROM2[221]<=26'd11274496; ROM3[221]<=26'd9735537; ROM4[221]<=26'd23442600;
ROM1[222]<=26'd1921798; ROM2[222]<=26'd11277983; ROM3[222]<=26'd9740933; ROM4[222]<=26'd23445207;
ROM1[223]<=26'd1932007; ROM2[223]<=26'd11284909; ROM3[223]<=26'd9745947; ROM4[223]<=26'd23451259;
ROM1[224]<=26'd1940249; ROM2[224]<=26'd11283735; ROM3[224]<=26'd9741833; ROM4[224]<=26'd23449158;
ROM1[225]<=26'd1947619; ROM2[225]<=26'd11283883; ROM3[225]<=26'd9734984; ROM4[225]<=26'd23445971;
ROM1[226]<=26'd1949077; ROM2[226]<=26'd11286577; ROM3[226]<=26'd9737211; ROM4[226]<=26'd23448139;
ROM1[227]<=26'd1941795; ROM2[227]<=26'd11285794; ROM3[227]<=26'd9738413; ROM4[227]<=26'd23447738;
ROM1[228]<=26'd1938949; ROM2[228]<=26'd11289185; ROM3[228]<=26'd9744764; ROM4[228]<=26'd23451784;
ROM1[229]<=26'd1936287; ROM2[229]<=26'd11291879; ROM3[229]<=26'd9749359; ROM4[229]<=26'd23454925;
ROM1[230]<=26'd1920800; ROM2[230]<=26'd11283790; ROM3[230]<=26'd9742094; ROM4[230]<=26'd23446394;
ROM1[231]<=26'd1917656; ROM2[231]<=26'd11279578; ROM3[231]<=26'd9735698; ROM4[231]<=26'd23441416;
ROM1[232]<=26'd1924418; ROM2[232]<=26'd11278667; ROM3[232]<=26'd9728968; ROM4[232]<=26'd23438873;
ROM1[233]<=26'd1936592; ROM2[233]<=26'd11278476; ROM3[233]<=26'd9723268; ROM4[233]<=26'd23437283;
ROM1[234]<=26'd1944026; ROM2[234]<=26'd11282768; ROM3[234]<=26'd9724789; ROM4[234]<=26'd23440779;
ROM1[235]<=26'd1939714; ROM2[235]<=26'd11284694; ROM3[235]<=26'd9728038; ROM4[235]<=26'd23441749;
ROM1[236]<=26'd1930657; ROM2[236]<=26'd11283270; ROM3[236]<=26'd9730959; ROM4[236]<=26'd23441600;
ROM1[237]<=26'd1924034; ROM2[237]<=26'd11281416; ROM3[237]<=26'd9732048; ROM4[237]<=26'd23441314;
ROM1[238]<=26'd1920664; ROM2[238]<=26'd11282716; ROM3[238]<=26'd9735511; ROM4[238]<=26'd23443395;
ROM1[239]<=26'd1921386; ROM2[239]<=26'd11285160; ROM3[239]<=26'd9739855; ROM4[239]<=26'd23446837;
ROM1[240]<=26'd1923880; ROM2[240]<=26'd11283562; ROM3[240]<=26'd9734367; ROM4[240]<=26'd23442994;
ROM1[241]<=26'd1938788; ROM2[241]<=26'd11285806; ROM3[241]<=26'd9730065; ROM4[241]<=26'd23443787;
ROM1[242]<=26'd1949930; ROM2[242]<=26'd11291193; ROM3[242]<=26'd9733336; ROM4[242]<=26'd23448098;
ROM1[243]<=26'd1934418; ROM2[243]<=26'd11280421; ROM3[243]<=26'd9726065; ROM4[243]<=26'd23439043;
ROM1[244]<=26'd1920368; ROM2[244]<=26'd11272431; ROM3[244]<=26'd9724190; ROM4[244]<=26'd23434483;
ROM1[245]<=26'd1917268; ROM2[245]<=26'd11274534; ROM3[245]<=26'd9730802; ROM4[245]<=26'd23438205;
ROM1[246]<=26'd1907587; ROM2[246]<=26'd11269222; ROM3[246]<=26'd9728102; ROM4[246]<=26'd23435440;
ROM1[247]<=26'd1910842; ROM2[247]<=26'd11274292; ROM3[247]<=26'd9733408; ROM4[247]<=26'd23439951;
ROM1[248]<=26'd1920952; ROM2[248]<=26'd11281169; ROM3[248]<=26'd9737748; ROM4[248]<=26'd23444701;
ROM1[249]<=26'd1926413; ROM2[249]<=26'd11281038; ROM3[249]<=26'd9731678; ROM4[249]<=26'd23440740;
ROM1[250]<=26'd1937271; ROM2[250]<=26'd11282585; ROM3[250]<=26'd9728726; ROM4[250]<=26'd23439226;
ROM1[251]<=26'd1933755; ROM2[251]<=26'd11281075; ROM3[251]<=26'd9727167; ROM4[251]<=26'd23438697;
ROM1[252]<=26'd1925528; ROM2[252]<=26'd11280509; ROM3[252]<=26'd9727848; ROM4[252]<=26'd23439081;
ROM1[253]<=26'd1921724; ROM2[253]<=26'd11281698; ROM3[253]<=26'd9732427; ROM4[253]<=26'd23439414;
ROM1[254]<=26'd1913091; ROM2[254]<=26'd11277588; ROM3[254]<=26'd9730300; ROM4[254]<=26'd23436512;
ROM1[255]<=26'd1906680; ROM2[255]<=26'd11274590; ROM3[255]<=26'd9730742; ROM4[255]<=26'd23436088;
ROM1[256]<=26'd1908871; ROM2[256]<=26'd11274782; ROM3[256]<=26'd9732256; ROM4[256]<=26'd23437792;
ROM1[257]<=26'd1914342; ROM2[257]<=26'd11270524; ROM3[257]<=26'd9724849; ROM4[257]<=26'd23436072;
ROM1[258]<=26'd1926385; ROM2[258]<=26'd11270219; ROM3[258]<=26'd9717422; ROM4[258]<=26'd23432548;
ROM1[259]<=26'd1933446; ROM2[259]<=26'd11275073; ROM3[259]<=26'd9717573; ROM4[259]<=26'd23433381;
ROM1[260]<=26'd1927778; ROM2[260]<=26'd11275490; ROM3[260]<=26'd9719594; ROM4[260]<=26'd23433414;
ROM1[261]<=26'd1920292; ROM2[261]<=26'd11275512; ROM3[261]<=26'd9723609; ROM4[261]<=26'd23433848;
ROM1[262]<=26'd1912947; ROM2[262]<=26'd11271397; ROM3[262]<=26'd9726362; ROM4[262]<=26'd23434985;
ROM1[263]<=26'd1903725; ROM2[263]<=26'd11267478; ROM3[263]<=26'd9728135; ROM4[263]<=26'd23432657;
ROM1[264]<=26'd1904705; ROM2[264]<=26'd11270487; ROM3[264]<=26'd9732312; ROM4[264]<=26'd23435289;
ROM1[265]<=26'd1914543; ROM2[265]<=26'd11275367; ROM3[265]<=26'd9733607; ROM4[265]<=26'd23438403;
ROM1[266]<=26'd1931749; ROM2[266]<=26'd11282603; ROM3[266]<=26'd9733145; ROM4[266]<=26'd23442754;
ROM1[267]<=26'd1946445; ROM2[267]<=26'd11290404; ROM3[267]<=26'd9736960; ROM4[267]<=26'd23450581;
ROM1[268]<=26'd1947128; ROM2[268]<=26'd11292333; ROM3[268]<=26'd9741976; ROM4[268]<=26'd23453928;
ROM1[269]<=26'd1937174; ROM2[269]<=26'd11287102; ROM3[269]<=26'd9740475; ROM4[269]<=26'd23451696;
ROM1[270]<=26'd1928970; ROM2[270]<=26'd11285172; ROM3[270]<=26'd9739804; ROM4[270]<=26'd23449176;
ROM1[271]<=26'd1921094; ROM2[271]<=26'd11282983; ROM3[271]<=26'd9742250; ROM4[271]<=26'd23447304;
ROM1[272]<=26'd1914936; ROM2[272]<=26'd11278991; ROM3[272]<=26'd9739669; ROM4[272]<=26'd23444487;
ROM1[273]<=26'd1919621; ROM2[273]<=26'd11280187; ROM3[273]<=26'd9739344; ROM4[273]<=26'd23445005;
ROM1[274]<=26'd1932397; ROM2[274]<=26'd11282741; ROM3[274]<=26'd9737219; ROM4[274]<=26'd23447010;
ROM1[275]<=26'd1939533; ROM2[275]<=26'd11280278; ROM3[275]<=26'd9727409; ROM4[275]<=26'd23442642;
ROM1[276]<=26'd1936294; ROM2[276]<=26'd11278580; ROM3[276]<=26'd9726065; ROM4[276]<=26'd23440542;
ROM1[277]<=26'd1934074; ROM2[277]<=26'd11281135; ROM3[277]<=26'd9732860; ROM4[277]<=26'd23443575;
ROM1[278]<=26'd1928921; ROM2[278]<=26'd11281826; ROM3[278]<=26'd9737386; ROM4[278]<=26'd23445059;
ROM1[279]<=26'd1930943; ROM2[279]<=26'd11287418; ROM3[279]<=26'd9744202; ROM4[279]<=26'd23450898;
ROM1[280]<=26'd1927186; ROM2[280]<=26'd11287377; ROM3[280]<=26'd9745601; ROM4[280]<=26'd23449509;
ROM1[281]<=26'd1920892; ROM2[281]<=26'd11283640; ROM3[281]<=26'd9740746; ROM4[281]<=26'd23444304;
ROM1[282]<=26'd1929105; ROM2[282]<=26'd11284447; ROM3[282]<=26'd9736718; ROM4[282]<=26'd23442848;
ROM1[283]<=26'd1936802; ROM2[283]<=26'd11280399; ROM3[283]<=26'd9728664; ROM4[283]<=26'd23439538;
ROM1[284]<=26'd1933948; ROM2[284]<=26'd11277634; ROM3[284]<=26'd9726403; ROM4[284]<=26'd23438089;
ROM1[285]<=26'd1927708; ROM2[285]<=26'd11277361; ROM3[285]<=26'd9727563; ROM4[285]<=26'd23437016;
ROM1[286]<=26'd1923577; ROM2[286]<=26'd11279389; ROM3[286]<=26'd9733161; ROM4[286]<=26'd23441392;
ROM1[287]<=26'd1921882; ROM2[287]<=26'd11283065; ROM3[287]<=26'd9740565; ROM4[287]<=26'd23446323;
ROM1[288]<=26'd1915573; ROM2[288]<=26'd11282210; ROM3[288]<=26'd9740571; ROM4[288]<=26'd23444736;
ROM1[289]<=26'd1909442; ROM2[289]<=26'd11275757; ROM3[289]<=26'd9735690; ROM4[289]<=26'd23439514;
ROM1[290]<=26'd1912493; ROM2[290]<=26'd11271600; ROM3[290]<=26'd9730635; ROM4[290]<=26'd23435931;
ROM1[291]<=26'd1924245; ROM2[291]<=26'd11273216; ROM3[291]<=26'd9726013; ROM4[291]<=26'd23436648;
ROM1[292]<=26'd1936227; ROM2[292]<=26'd11276539; ROM3[292]<=26'd9725963; ROM4[292]<=26'd23440920;
ROM1[293]<=26'd1938124; ROM2[293]<=26'd11281800; ROM3[293]<=26'd9733122; ROM4[293]<=26'd23446000;
ROM1[294]<=26'd1934287; ROM2[294]<=26'd11287149; ROM3[294]<=26'd9741428; ROM4[294]<=26'd23449400;
ROM1[295]<=26'd1928458; ROM2[295]<=26'd11286830; ROM3[295]<=26'd9743851; ROM4[295]<=26'd23449536;
ROM1[296]<=26'd1922777; ROM2[296]<=26'd11286380; ROM3[296]<=26'd9745086; ROM4[296]<=26'd23451138;
ROM1[297]<=26'd1912841; ROM2[297]<=26'd11278872; ROM3[297]<=26'd9739160; ROM4[297]<=26'd23443340;
ROM1[298]<=26'd1907962; ROM2[298]<=26'd11269659; ROM3[298]<=26'd9728437; ROM4[298]<=26'd23434445;
ROM1[299]<=26'd1918460; ROM2[299]<=26'd11271777; ROM3[299]<=26'd9723005; ROM4[299]<=26'd23434386;
ROM1[300]<=26'd1926833; ROM2[300]<=26'd11272583; ROM3[300]<=26'd9718108; ROM4[300]<=26'd23433298;
ROM1[301]<=26'd1927135; ROM2[301]<=26'd11274929; ROM3[301]<=26'd9720941; ROM4[301]<=26'd23437287;
ROM1[302]<=26'd1918454; ROM2[302]<=26'd11274282; ROM3[302]<=26'd9723180; ROM4[302]<=26'd23436565;
ROM1[303]<=26'd1909752; ROM2[303]<=26'd11270918; ROM3[303]<=26'd9725453; ROM4[303]<=26'd23435106;
ROM1[304]<=26'd1909412; ROM2[304]<=26'd11274174; ROM3[304]<=26'd9731958; ROM4[304]<=26'd23437910;
ROM1[305]<=26'd1910942; ROM2[305]<=26'd11279717; ROM3[305]<=26'd9738804; ROM4[305]<=26'd23442421;
ROM1[306]<=26'd1913917; ROM2[306]<=26'd11281723; ROM3[306]<=26'd9742027; ROM4[306]<=26'd23445007;
ROM1[307]<=26'd1919615; ROM2[307]<=26'd11278370; ROM3[307]<=26'd9734781; ROM4[307]<=26'd23440446;
ROM1[308]<=26'd1931623; ROM2[308]<=26'd11278421; ROM3[308]<=26'd9726471; ROM4[308]<=26'd23437707;
ROM1[309]<=26'd1932461; ROM2[309]<=26'd11276353; ROM3[309]<=26'd9723223; ROM4[309]<=26'd23436145;
ROM1[310]<=26'd1926029; ROM2[310]<=26'd11275425; ROM3[310]<=26'd9725621; ROM4[310]<=26'd23437373;
ROM1[311]<=26'd1923373; ROM2[311]<=26'd11280507; ROM3[311]<=26'd9732602; ROM4[311]<=26'd23441093;
ROM1[312]<=26'd1922919; ROM2[312]<=26'd11284731; ROM3[312]<=26'd9739610; ROM4[312]<=26'd23445299;
ROM1[313]<=26'd1924211; ROM2[313]<=26'd11291868; ROM3[313]<=26'd9749433; ROM4[313]<=26'd23452936;
ROM1[314]<=26'd1926640; ROM2[314]<=26'd11292677; ROM3[314]<=26'd9750311; ROM4[314]<=26'd23453145;
ROM1[315]<=26'd1925797; ROM2[315]<=26'd11285421; ROM3[315]<=26'd9741736; ROM4[315]<=26'd23446350;
ROM1[316]<=26'd1937341; ROM2[316]<=26'd11285768; ROM3[316]<=26'd9737270; ROM4[316]<=26'd23445302;
ROM1[317]<=26'd1945922; ROM2[317]<=26'd11286757; ROM3[317]<=26'd9731859; ROM4[317]<=26'd23444401;
ROM1[318]<=26'd1938802; ROM2[318]<=26'd11284541; ROM3[318]<=26'd9728552; ROM4[318]<=26'd23441447;
ROM1[319]<=26'd1930891; ROM2[319]<=26'd11284591; ROM3[319]<=26'd9732216; ROM4[319]<=26'd23441190;
ROM1[320]<=26'd1925950; ROM2[320]<=26'd11286140; ROM3[320]<=26'd9736376; ROM4[320]<=26'd23444677;
ROM1[321]<=26'd1917521; ROM2[321]<=26'd11284335; ROM3[321]<=26'd9735803; ROM4[321]<=26'd23444005;
ROM1[322]<=26'd1913865; ROM2[322]<=26'd11284756; ROM3[322]<=26'd9737009; ROM4[322]<=26'd23444731;
ROM1[323]<=26'd1921820; ROM2[323]<=26'd11288216; ROM3[323]<=26'd9738480; ROM4[323]<=26'd23448171;
ROM1[324]<=26'd1930230; ROM2[324]<=26'd11287046; ROM3[324]<=26'd9731681; ROM4[324]<=26'd23444552;
ROM1[325]<=26'd1943286; ROM2[325]<=26'd11289134; ROM3[325]<=26'd9729797; ROM4[325]<=26'd23446226;
ROM1[326]<=26'd1949245; ROM2[326]<=26'd11293886; ROM3[326]<=26'd9735954; ROM4[326]<=26'd23452507;
ROM1[327]<=26'd1945394; ROM2[327]<=26'd11296705; ROM3[327]<=26'd9742189; ROM4[327]<=26'd23455286;
ROM1[328]<=26'd1930523; ROM2[328]<=26'd11287710; ROM3[328]<=26'd9740242; ROM4[328]<=26'd23448075;
ROM1[329]<=26'd1915290; ROM2[329]<=26'd11277627; ROM3[329]<=26'd9735789; ROM4[329]<=26'd23439850;
ROM1[330]<=26'd1907238; ROM2[330]<=26'd11276837; ROM3[330]<=26'd9737205; ROM4[330]<=26'd23438925;
ROM1[331]<=26'd1911713; ROM2[331]<=26'd11277965; ROM3[331]<=26'd9738963; ROM4[331]<=26'd23440741;
ROM1[332]<=26'd1927703; ROM2[332]<=26'd11282962; ROM3[332]<=26'd9740558; ROM4[332]<=26'd23445081;
ROM1[333]<=26'd1944035; ROM2[333]<=26'd11288803; ROM3[333]<=26'd9740875; ROM4[333]<=26'd23450006;
ROM1[334]<=26'd1949939; ROM2[334]<=26'd11291066; ROM3[334]<=26'd9743256; ROM4[334]<=26'd23451220;
ROM1[335]<=26'd1937545; ROM2[335]<=26'd11283964; ROM3[335]<=26'd9738723; ROM4[335]<=26'd23446105;
ROM1[336]<=26'd1924250; ROM2[336]<=26'd11277989; ROM3[336]<=26'd9736987; ROM4[336]<=26'd23443600;
ROM1[337]<=26'd1920715; ROM2[337]<=26'd11279398; ROM3[337]<=26'd9740644; ROM4[337]<=26'd23444189;
ROM1[338]<=26'd1914327; ROM2[338]<=26'd11277306; ROM3[338]<=26'd9740684; ROM4[338]<=26'd23442425;
ROM1[339]<=26'd1913380; ROM2[339]<=26'd11277872; ROM3[339]<=26'd9743698; ROM4[339]<=26'd23443681;
ROM1[340]<=26'd1921232; ROM2[340]<=26'd11280176; ROM3[340]<=26'd9743424; ROM4[340]<=26'd23444800;
ROM1[341]<=26'd1933148; ROM2[341]<=26'd11280604; ROM3[341]<=26'd9735264; ROM4[341]<=26'd23443104;
ROM1[342]<=26'd1934624; ROM2[342]<=26'd11274512; ROM3[342]<=26'd9725805; ROM4[342]<=26'd23437500;
ROM1[343]<=26'd1930068; ROM2[343]<=26'd11271587; ROM3[343]<=26'd9724911; ROM4[343]<=26'd23434496;
ROM1[344]<=26'd1924550; ROM2[344]<=26'd11273442; ROM3[344]<=26'd9728414; ROM4[344]<=26'd23436508;
ROM1[345]<=26'd1918034; ROM2[345]<=26'd11272951; ROM3[345]<=26'd9730911; ROM4[345]<=26'd23437101;
ROM1[346]<=26'd1913110; ROM2[346]<=26'd11274503; ROM3[346]<=26'd9734862; ROM4[346]<=26'd23438811;
ROM1[347]<=26'd1912761; ROM2[347]<=26'd11277563; ROM3[347]<=26'd9738126; ROM4[347]<=26'd23441836;
ROM1[348]<=26'd1915612; ROM2[348]<=26'd11277503; ROM3[348]<=26'd9735009; ROM4[348]<=26'd23439904;
ROM1[349]<=26'd1925954; ROM2[349]<=26'd11276516; ROM3[349]<=26'd9730278; ROM4[349]<=26'd23439555;
ROM1[350]<=26'd1938707; ROM2[350]<=26'd11278522; ROM3[350]<=26'd9728173; ROM4[350]<=26'd23442061;
ROM1[351]<=26'd1940327; ROM2[351]<=26'd11281134; ROM3[351]<=26'd9731843; ROM4[351]<=26'd23445155;
ROM1[352]<=26'd1936709; ROM2[352]<=26'd11281677; ROM3[352]<=26'd9738858; ROM4[352]<=26'd23448773;
ROM1[353]<=26'd1927962; ROM2[353]<=26'd11279566; ROM3[353]<=26'd9742261; ROM4[353]<=26'd23447368;
ROM1[354]<=26'd1921781; ROM2[354]<=26'd11279355; ROM3[354]<=26'd9743507; ROM4[354]<=26'd23446592;
ROM1[355]<=26'd1916309; ROM2[355]<=26'd11278075; ROM3[355]<=26'd9743629; ROM4[355]<=26'd23445194;
ROM1[356]<=26'd1916083; ROM2[356]<=26'd11276336; ROM3[356]<=26'd9742139; ROM4[356]<=26'd23443626;
ROM1[357]<=26'd1924859; ROM2[357]<=26'd11277921; ROM3[357]<=26'd9738882; ROM4[357]<=26'd23444985;
ROM1[358]<=26'd1937988; ROM2[358]<=26'd11280939; ROM3[358]<=26'd9733859; ROM4[358]<=26'd23446741;
ROM1[359]<=26'd1937343; ROM2[359]<=26'd11278748; ROM3[359]<=26'd9729596; ROM4[359]<=26'd23444065;
ROM1[360]<=26'd1929281; ROM2[360]<=26'd11276841; ROM3[360]<=26'd9729512; ROM4[360]<=26'd23442099;
ROM1[361]<=26'd1927284; ROM2[361]<=26'd11282236; ROM3[361]<=26'd9737755; ROM4[361]<=26'd23447070;
ROM1[362]<=26'd1930412; ROM2[362]<=26'd11290108; ROM3[362]<=26'd9748383; ROM4[362]<=26'd23454999;
ROM1[363]<=26'd1918710; ROM2[363]<=26'd11283738; ROM3[363]<=26'd9745125; ROM4[363]<=26'd23452016;
ROM1[364]<=26'd1912427; ROM2[364]<=26'd11278456; ROM3[364]<=26'd9741491; ROM4[364]<=26'd23447939;
ROM1[365]<=26'd1921304; ROM2[365]<=26'd11279679; ROM3[365]<=26'd9739718; ROM4[365]<=26'd23447373;
ROM1[366]<=26'd1931931; ROM2[366]<=26'd11278234; ROM3[366]<=26'd9731413; ROM4[366]<=26'd23443408;
ROM1[367]<=26'd1947657; ROM2[367]<=26'd11286218; ROM3[367]<=26'd9734737; ROM4[367]<=26'd23449666;
ROM1[368]<=26'd1953174; ROM2[368]<=26'd11293879; ROM3[368]<=26'd9743728; ROM4[368]<=26'd23457334;
ROM1[369]<=26'd1943246; ROM2[369]<=26'd11292269; ROM3[369]<=26'd9744807; ROM4[369]<=26'd23456216;
ROM1[370]<=26'd1932096; ROM2[370]<=26'd11287618; ROM3[370]<=26'd9745324; ROM4[370]<=26'd23452875;
ROM1[371]<=26'd1919512; ROM2[371]<=26'd11281678; ROM3[371]<=26'd9742696; ROM4[371]<=26'd23447129;
ROM1[372]<=26'd1916016; ROM2[372]<=26'd11282090; ROM3[372]<=26'd9741244; ROM4[372]<=26'd23444975;
ROM1[373]<=26'd1920981; ROM2[373]<=26'd11283085; ROM3[373]<=26'd9738425; ROM4[373]<=26'd23442395;
ROM1[374]<=26'd1930604; ROM2[374]<=26'd11282481; ROM3[374]<=26'd9733381; ROM4[374]<=26'd23441222;
ROM1[375]<=26'd1944073; ROM2[375]<=26'd11286401; ROM3[375]<=26'd9735450; ROM4[375]<=26'd23446408;
ROM1[376]<=26'd1942222; ROM2[376]<=26'd11285825; ROM3[376]<=26'd9738480; ROM4[376]<=26'd23447858;
ROM1[377]<=26'd1933404; ROM2[377]<=26'd11281909; ROM3[377]<=26'd9739989; ROM4[377]<=26'd23446064;
ROM1[378]<=26'd1927250; ROM2[378]<=26'd11279916; ROM3[378]<=26'd9740964; ROM4[378]<=26'd23444391;
ROM1[379]<=26'd1921955; ROM2[379]<=26'd11281881; ROM3[379]<=26'd9742919; ROM4[379]<=26'd23444713;
ROM1[380]<=26'd1918534; ROM2[380]<=26'd11284627; ROM3[380]<=26'd9745742; ROM4[380]<=26'd23446444;
ROM1[381]<=26'd1922894; ROM2[381]<=26'd11287754; ROM3[381]<=26'd9750682; ROM4[381]<=26'd23450752;
ROM1[382]<=26'd1939949; ROM2[382]<=26'd11296412; ROM3[382]<=26'd9755988; ROM4[382]<=26'd23459216;
ROM1[383]<=26'd1954221; ROM2[383]<=26'd11298942; ROM3[383]<=26'd9749932; ROM4[383]<=26'd23458806;
ROM1[384]<=26'd1945612; ROM2[384]<=26'd11286509; ROM3[384]<=26'd9735823; ROM4[384]<=26'd23446448;
ROM1[385]<=26'd1933624; ROM2[385]<=26'd11279707; ROM3[385]<=26'd9733460; ROM4[385]<=26'd23441742;
ROM1[386]<=26'd1927125; ROM2[386]<=26'd11282575; ROM3[386]<=26'd9738002; ROM4[386]<=26'd23443206;
ROM1[387]<=26'd1922224; ROM2[387]<=26'd11280655; ROM3[387]<=26'd9740200; ROM4[387]<=26'd23441517;
ROM1[388]<=26'd1916598; ROM2[388]<=26'd11279999; ROM3[388]<=26'd9743335; ROM4[388]<=26'd23442597;
ROM1[389]<=26'd1914623; ROM2[389]<=26'd11280532; ROM3[389]<=26'd9740664; ROM4[389]<=26'd23440302;
ROM1[390]<=26'd1915164; ROM2[390]<=26'd11274837; ROM3[390]<=26'd9733836; ROM4[390]<=26'd23433221;
ROM1[391]<=26'd1929653; ROM2[391]<=26'd11277271; ROM3[391]<=26'd9729189; ROM4[391]<=26'd23433752;
ROM1[392]<=26'd1942660; ROM2[392]<=26'd11283115; ROM3[392]<=26'd9730795; ROM4[392]<=26'd23439353;
ROM1[393]<=26'd1937768; ROM2[393]<=26'd11282068; ROM3[393]<=26'd9731968; ROM4[393]<=26'd23439480;
ROM1[394]<=26'd1927283; ROM2[394]<=26'd11277583; ROM3[394]<=26'd9730321; ROM4[394]<=26'd23435261;
ROM1[395]<=26'd1922239; ROM2[395]<=26'd11276782; ROM3[395]<=26'd9734241; ROM4[395]<=26'd23436679;
ROM1[396]<=26'd1917837; ROM2[396]<=26'd11277300; ROM3[396]<=26'd9736977; ROM4[396]<=26'd23437401;
ROM1[397]<=26'd1915574; ROM2[397]<=26'd11277220; ROM3[397]<=26'd9737710; ROM4[397]<=26'd23436417;
ROM1[398]<=26'd1922575; ROM2[398]<=26'd11281669; ROM3[398]<=26'd9740349; ROM4[398]<=26'd23441220;
ROM1[399]<=26'd1934645; ROM2[399]<=26'd11285922; ROM3[399]<=26'd9735775; ROM4[399]<=26'd23441823;
ROM1[400]<=26'd1944703; ROM2[400]<=26'd11287373; ROM3[400]<=26'd9728395; ROM4[400]<=26'd23439840;
ROM1[401]<=26'd1941002; ROM2[401]<=26'd11283870; ROM3[401]<=26'd9726948; ROM4[401]<=26'd23437705;
ROM1[402]<=26'd1930670; ROM2[402]<=26'd11279628; ROM3[402]<=26'd9726491; ROM4[402]<=26'd23435251;
ROM1[403]<=26'd1924168; ROM2[403]<=26'd11279588; ROM3[403]<=26'd9730879; ROM4[403]<=26'd23436394;
ROM1[404]<=26'd1918705; ROM2[404]<=26'd11280068; ROM3[404]<=26'd9738470; ROM4[404]<=26'd23440094;
ROM1[405]<=26'd1915822; ROM2[405]<=26'd11282033; ROM3[405]<=26'd9742547; ROM4[405]<=26'd23443417;
ROM1[406]<=26'd1919237; ROM2[406]<=26'd11283191; ROM3[406]<=26'd9742683; ROM4[406]<=26'd23444109;
ROM1[407]<=26'd1928141; ROM2[407]<=26'd11283576; ROM3[407]<=26'd9740544; ROM4[407]<=26'd23445570;
ROM1[408]<=26'd1941541; ROM2[408]<=26'd11284364; ROM3[408]<=26'd9736036; ROM4[408]<=26'd23445470;
ROM1[409]<=26'd1953282; ROM2[409]<=26'd11291104; ROM3[409]<=26'd9743279; ROM4[409]<=26'd23453513;
ROM1[410]<=26'd1952597; ROM2[410]<=26'd11294315; ROM3[410]<=26'd9750956; ROM4[410]<=26'd23459211;
ROM1[411]<=26'd1938276; ROM2[411]<=26'd11285569; ROM3[411]<=26'd9747158; ROM4[411]<=26'd23451974;
ROM1[412]<=26'd1936219; ROM2[412]<=26'd11286624; ROM3[412]<=26'd9751645; ROM4[412]<=26'd23455591;
ROM1[413]<=26'd1929172; ROM2[413]<=26'd11284567; ROM3[413]<=26'd9753700; ROM4[413]<=26'd23455650;
ROM1[414]<=26'd1925360; ROM2[414]<=26'd11281211; ROM3[414]<=26'd9752249; ROM4[414]<=26'd23453909;
ROM1[415]<=26'd1936986; ROM2[415]<=26'd11286878; ROM3[415]<=26'd9752895; ROM4[415]<=26'd23457821;
ROM1[416]<=26'd1950690; ROM2[416]<=26'd11287576; ROM3[416]<=26'd9747790; ROM4[416]<=26'd23455781;
ROM1[417]<=26'd1955409; ROM2[417]<=26'd11286814; ROM3[417]<=26'd9743041; ROM4[417]<=26'd23455442;
ROM1[418]<=26'd1953597; ROM2[418]<=26'd11290157; ROM3[418]<=26'd9749636; ROM4[418]<=26'd23460300;
ROM1[419]<=26'd1947396; ROM2[419]<=26'd11291491; ROM3[419]<=26'd9755131; ROM4[419]<=26'd23462021;
ROM1[420]<=26'd1936237; ROM2[420]<=26'd11288227; ROM3[420]<=26'd9752755; ROM4[420]<=26'd23457288;
ROM1[421]<=26'd1927670; ROM2[421]<=26'd11284748; ROM3[421]<=26'd9751549; ROM4[421]<=26'd23453340;
ROM1[422]<=26'd1921533; ROM2[422]<=26'd11280591; ROM3[422]<=26'd9747200; ROM4[422]<=26'd23448560;
ROM1[423]<=26'd1927930; ROM2[423]<=26'd11282022; ROM3[423]<=26'd9747668; ROM4[423]<=26'd23450424;
ROM1[424]<=26'd1940397; ROM2[424]<=26'd11285977; ROM3[424]<=26'd9746511; ROM4[424]<=26'd23453867;
ROM1[425]<=26'd1945183; ROM2[425]<=26'd11283021; ROM3[425]<=26'd9738964; ROM4[425]<=26'd23450290;
ROM1[426]<=26'd1943736; ROM2[426]<=26'd11281868; ROM3[426]<=26'd9738351; ROM4[426]<=26'd23449243;
ROM1[427]<=26'd1936903; ROM2[427]<=26'd11282525; ROM3[427]<=26'd9742716; ROM4[427]<=26'd23450043;
ROM1[428]<=26'd1930709; ROM2[428]<=26'd11281966; ROM3[428]<=26'd9747680; ROM4[428]<=26'd23451357;
ROM1[429]<=26'd1929634; ROM2[429]<=26'd11284096; ROM3[429]<=26'd9753414; ROM4[429]<=26'd23455318;
ROM1[430]<=26'd1929073; ROM2[430]<=26'd11286917; ROM3[430]<=26'd9758390; ROM4[430]<=26'd23458769;
ROM1[431]<=26'd1931436; ROM2[431]<=26'd11285739; ROM3[431]<=26'd9759932; ROM4[431]<=26'd23460014;
ROM1[432]<=26'd1943701; ROM2[432]<=26'd11288003; ROM3[432]<=26'd9760642; ROM4[432]<=26'd23462271;
ROM1[433]<=26'd1957501; ROM2[433]<=26'd11291597; ROM3[433]<=26'd9757489; ROM4[433]<=26'd23462579;
ROM1[434]<=26'd1946284; ROM2[434]<=26'd11277726; ROM3[434]<=26'd9743626; ROM4[434]<=26'd23450995;
ROM1[435]<=26'd1931119; ROM2[435]<=26'd11267531; ROM3[435]<=26'd9737029; ROM4[435]<=26'd23443501;
ROM1[436]<=26'd1926336; ROM2[436]<=26'd11269452; ROM3[436]<=26'd9740948; ROM4[436]<=26'd23444910;
ROM1[437]<=26'd1924611; ROM2[437]<=26'd11272407; ROM3[437]<=26'd9744609; ROM4[437]<=26'd23446649;
ROM1[438]<=26'd1923853; ROM2[438]<=26'd11277998; ROM3[438]<=26'd9752624; ROM4[438]<=26'd23452194;
ROM1[439]<=26'd1925754; ROM2[439]<=26'd11280622; ROM3[439]<=26'd9755116; ROM4[439]<=26'd23454141;
ROM1[440]<=26'd1936936; ROM2[440]<=26'd11284961; ROM3[440]<=26'd9754884; ROM4[440]<=26'd23456330;
ROM1[441]<=26'd1956220; ROM2[441]<=26'd11292783; ROM3[441]<=26'd9757881; ROM4[441]<=26'd23464163;
ROM1[442]<=26'd1966128; ROM2[442]<=26'd11296788; ROM3[442]<=26'd9760068; ROM4[442]<=26'd23467296;
ROM1[443]<=26'd1957483; ROM2[443]<=26'd11291957; ROM3[443]<=26'd9758083; ROM4[443]<=26'd23463440;
ROM1[444]<=26'd1943208; ROM2[444]<=26'd11282568; ROM3[444]<=26'd9754271; ROM4[444]<=26'd23455845;
ROM1[445]<=26'd1933298; ROM2[445]<=26'd11274849; ROM3[445]<=26'd9749946; ROM4[445]<=26'd23450717;
ROM1[446]<=26'd1926305; ROM2[446]<=26'd11272144; ROM3[446]<=26'd9750731; ROM4[446]<=26'd23449221;
ROM1[447]<=26'd1926167; ROM2[447]<=26'd11276917; ROM3[447]<=26'd9757102; ROM4[447]<=26'd23452027;
ROM1[448]<=26'd1926453; ROM2[448]<=26'd11277860; ROM3[448]<=26'd9754546; ROM4[448]<=26'd23451773;
ROM1[449]<=26'd1934628; ROM2[449]<=26'd11276861; ROM3[449]<=26'd9747306; ROM4[449]<=26'd23448376;
ROM1[450]<=26'd1946846; ROM2[450]<=26'd11279222; ROM3[450]<=26'd9742795; ROM4[450]<=26'd23448084;
ROM1[451]<=26'd1944298; ROM2[451]<=26'd11278109; ROM3[451]<=26'd9740576; ROM4[451]<=26'd23446760;
ROM1[452]<=26'd1940481; ROM2[452]<=26'd11280642; ROM3[452]<=26'd9745892; ROM4[452]<=26'd23450072;
ROM1[453]<=26'd1938095; ROM2[453]<=26'd11283336; ROM3[453]<=26'd9751906; ROM4[453]<=26'd23452232;
ROM1[454]<=26'd1932201; ROM2[454]<=26'd11282185; ROM3[454]<=26'd9752149; ROM4[454]<=26'd23450503;
ROM1[455]<=26'd1927500; ROM2[455]<=26'd11282583; ROM3[455]<=26'd9754857; ROM4[455]<=26'd23449965;
ROM1[456]<=26'd1928808; ROM2[456]<=26'd11281134; ROM3[456]<=26'd9753193; ROM4[456]<=26'd23448376;
ROM1[457]<=26'd1934232; ROM2[457]<=26'd11278224; ROM3[457]<=26'd9744667; ROM4[457]<=26'd23444678;
ROM1[458]<=26'd1947974; ROM2[458]<=26'd11280817; ROM3[458]<=26'd9740956; ROM4[458]<=26'd23446464;
ROM1[459]<=26'd1953977; ROM2[459]<=26'd11283234; ROM3[459]<=26'd9741438; ROM4[459]<=26'd23450419;
ROM1[460]<=26'd1946889; ROM2[460]<=26'd11281190; ROM3[460]<=26'd9744228; ROM4[460]<=26'd23451448;
ROM1[461]<=26'd1939397; ROM2[461]<=26'd11280078; ROM3[461]<=26'd9748202; ROM4[461]<=26'd23451297;
ROM1[462]<=26'd1932166; ROM2[462]<=26'd11276734; ROM3[462]<=26'd9748532; ROM4[462]<=26'd23449006;
ROM1[463]<=26'd1926575; ROM2[463]<=26'd11276836; ROM3[463]<=26'd9751907; ROM4[463]<=26'd23449168;
ROM1[464]<=26'd1925742; ROM2[464]<=26'd11279583; ROM3[464]<=26'd9753294; ROM4[464]<=26'd23450296;
ROM1[465]<=26'd1929208; ROM2[465]<=26'd11279268; ROM3[465]<=26'd9749076; ROM4[465]<=26'd23450024;
ROM1[466]<=26'd1943341; ROM2[466]<=26'd11281033; ROM3[466]<=26'd9746562; ROM4[466]<=26'd23451987;
ROM1[467]<=26'd1953149; ROM2[467]<=26'd11283026; ROM3[467]<=26'd9745570; ROM4[467]<=26'd23453181;
ROM1[468]<=26'd1945213; ROM2[468]<=26'd11278514; ROM3[468]<=26'd9741286; ROM4[468]<=26'd23448106;
ROM1[469]<=26'd1941158; ROM2[469]<=26'd11279969; ROM3[469]<=26'd9746492; ROM4[469]<=26'd23449489;
ROM1[470]<=26'd1939272; ROM2[470]<=26'd11283631; ROM3[470]<=26'd9751210; ROM4[470]<=26'd23452597;
ROM1[471]<=26'd1931523; ROM2[471]<=26'd11281424; ROM3[471]<=26'd9750076; ROM4[471]<=26'd23451895;
ROM1[472]<=26'd1928128; ROM2[472]<=26'd11280903; ROM3[472]<=26'd9751023; ROM4[472]<=26'd23451774;
ROM1[473]<=26'd1927970; ROM2[473]<=26'd11277237; ROM3[473]<=26'd9748824; ROM4[473]<=26'd23448821;
ROM1[474]<=26'd1936794; ROM2[474]<=26'd11274530; ROM3[474]<=26'd9745530; ROM4[474]<=26'd23445216;
ROM1[475]<=26'd1947203; ROM2[475]<=26'd11274513; ROM3[475]<=26'd9742008; ROM4[475]<=26'd23444186;
ROM1[476]<=26'd1949899; ROM2[476]<=26'd11277957; ROM3[476]<=26'd9746465; ROM4[476]<=26'd23447240;
ROM1[477]<=26'd1948799; ROM2[477]<=26'd11284123; ROM3[477]<=26'd9756494; ROM4[477]<=26'd23454727;
ROM1[478]<=26'd1938330; ROM2[478]<=26'd11280676; ROM3[478]<=26'd9757690; ROM4[478]<=26'd23453842;
ROM1[479]<=26'd1926098; ROM2[479]<=26'd11272554; ROM3[479]<=26'd9754720; ROM4[479]<=26'd23447406;
ROM1[480]<=26'd1926175; ROM2[480]<=26'd11275923; ROM3[480]<=26'd9761636; ROM4[480]<=26'd23452285;
ROM1[481]<=26'd1936432; ROM2[481]<=26'd11285462; ROM3[481]<=26'd9769245; ROM4[481]<=26'd23459989;
ROM1[482]<=26'd1940232; ROM2[482]<=26'd11282562; ROM3[482]<=26'd9758873; ROM4[482]<=26'd23453770;
ROM1[483]<=26'd1948005; ROM2[483]<=26'd11278865; ROM3[483]<=26'd9748011; ROM4[483]<=26'd23449173;
ROM1[484]<=26'd1946113; ROM2[484]<=26'd11273794; ROM3[484]<=26'd9742212; ROM4[484]<=26'd23445078;
ROM1[485]<=26'd1932685; ROM2[485]<=26'd11264705; ROM3[485]<=26'd9735959; ROM4[485]<=26'd23437871;
ROM1[486]<=26'd1927734; ROM2[486]<=26'd11265522; ROM3[486]<=26'd9740363; ROM4[486]<=26'd23440350;
ROM1[487]<=26'd1927175; ROM2[487]<=26'd11271754; ROM3[487]<=26'd9747633; ROM4[487]<=26'd23444301;
ROM1[488]<=26'd1921121; ROM2[488]<=26'd11272588; ROM3[488]<=26'd9749897; ROM4[488]<=26'd23444992;
ROM1[489]<=26'd1920141; ROM2[489]<=26'd11271809; ROM3[489]<=26'd9747355; ROM4[489]<=26'd23442984;
ROM1[490]<=26'd1929186; ROM2[490]<=26'd11277930; ROM3[490]<=26'd9746897; ROM4[490]<=26'd23445588;
ROM1[491]<=26'd1940712; ROM2[491]<=26'd11280650; ROM3[491]<=26'd9741804; ROM4[491]<=26'd23446469;
ROM1[492]<=26'd1946470; ROM2[492]<=26'd11279045; ROM3[492]<=26'd9737837; ROM4[492]<=26'd23444962;
ROM1[493]<=26'd1940002; ROM2[493]<=26'd11277304; ROM3[493]<=26'd9737335; ROM4[493]<=26'd23444599;
ROM1[494]<=26'd1931912; ROM2[494]<=26'd11277444; ROM3[494]<=26'd9740782; ROM4[494]<=26'd23445944;
ROM1[495]<=26'd1927365; ROM2[495]<=26'd11278810; ROM3[495]<=26'd9744714; ROM4[495]<=26'd23446909;
ROM1[496]<=26'd1923421; ROM2[496]<=26'd11279509; ROM3[496]<=26'd9748564; ROM4[496]<=26'd23449525;
ROM1[497]<=26'd1921301; ROM2[497]<=26'd11281616; ROM3[497]<=26'd9753121; ROM4[497]<=26'd23452027;
ROM1[498]<=26'd1925915; ROM2[498]<=26'd11282831; ROM3[498]<=26'd9751795; ROM4[498]<=26'd23451389;
ROM1[499]<=26'd1940011; ROM2[499]<=26'd11286089; ROM3[499]<=26'd9749556; ROM4[499]<=26'd23453792;
ROM1[500]<=26'd1954448; ROM2[500]<=26'd11292139; ROM3[500]<=26'd9747700; ROM4[500]<=26'd23457059;
ROM1[501]<=26'd1954345; ROM2[501]<=26'd11292801; ROM3[501]<=26'd9750053; ROM4[501]<=26'd23456783;
ROM1[502]<=26'd1946350; ROM2[502]<=26'd11289899; ROM3[502]<=26'd9751323; ROM4[502]<=26'd23455422;
ROM1[503]<=26'd1938515; ROM2[503]<=26'd11289521; ROM3[503]<=26'd9751021; ROM4[503]<=26'd23453288;
ROM1[504]<=26'd1932918; ROM2[504]<=26'd11289730; ROM3[504]<=26'd9752866; ROM4[504]<=26'd23452981;
ROM1[505]<=26'd1923426; ROM2[505]<=26'd11284447; ROM3[505]<=26'd9749665; ROM4[505]<=26'd23449032;
ROM1[506]<=26'd1923048; ROM2[506]<=26'd11281431; ROM3[506]<=26'd9747322; ROM4[506]<=26'd23445872;
ROM1[507]<=26'd1937583; ROM2[507]<=26'd11285080; ROM3[507]<=26'd9747981; ROM4[507]<=26'd23450663;
ROM1[508]<=26'd1951264; ROM2[508]<=26'd11284565; ROM3[508]<=26'd9744373; ROM4[508]<=26'd23451659;
ROM1[509]<=26'd1956946; ROM2[509]<=26'd11286685; ROM3[509]<=26'd9746618; ROM4[509]<=26'd23455234;
ROM1[510]<=26'd1954236; ROM2[510]<=26'd11290440; ROM3[510]<=26'd9752389; ROM4[510]<=26'd23458791;
ROM1[511]<=26'd1944810; ROM2[511]<=26'd11286920; ROM3[511]<=26'd9755068; ROM4[511]<=26'd23457720;
ROM1[512]<=26'd1935810; ROM2[512]<=26'd11283742; ROM3[512]<=26'd9755561; ROM4[512]<=26'd23454814;
ROM1[513]<=26'd1928139; ROM2[513]<=26'd11279453; ROM3[513]<=26'd9754950; ROM4[513]<=26'd23451386;
ROM1[514]<=26'd1932818; ROM2[514]<=26'd11284401; ROM3[514]<=26'd9761373; ROM4[514]<=26'd23458141;
ROM1[515]<=26'd1937832; ROM2[515]<=26'd11283998; ROM3[515]<=26'd9759067; ROM4[515]<=26'd23456822;
ROM1[516]<=26'd1942296; ROM2[516]<=26'd11278150; ROM3[516]<=26'd9747801; ROM4[516]<=26'd23449897;
ROM1[517]<=26'd1946981; ROM2[517]<=26'd11278977; ROM3[517]<=26'd9743294; ROM4[517]<=26'd23449038;
ROM1[518]<=26'd1940710; ROM2[518]<=26'd11276103; ROM3[518]<=26'd9740686; ROM4[518]<=26'd23446101;
ROM1[519]<=26'd1933563; ROM2[519]<=26'd11275278; ROM3[519]<=26'd9744825; ROM4[519]<=26'd23446061;
ROM1[520]<=26'd1931419; ROM2[520]<=26'd11277880; ROM3[520]<=26'd9751815; ROM4[520]<=26'd23449830;
ROM1[521]<=26'd1927061; ROM2[521]<=26'd11280317; ROM3[521]<=26'd9755560; ROM4[521]<=26'd23450159;
ROM1[522]<=26'd1928423; ROM2[522]<=26'd11284020; ROM3[522]<=26'd9759520; ROM4[522]<=26'd23455751;
ROM1[523]<=26'd1936427; ROM2[523]<=26'd11287410; ROM3[523]<=26'd9759999; ROM4[523]<=26'd23459880;
ROM1[524]<=26'd1943127; ROM2[524]<=26'd11284860; ROM3[524]<=26'd9752710; ROM4[524]<=26'd23454678;
ROM1[525]<=26'd1954182; ROM2[525]<=26'd11285561; ROM3[525]<=26'd9751100; ROM4[525]<=26'd23458759;
ROM1[526]<=26'd1947466; ROM2[526]<=26'd11278862; ROM3[526]<=26'd9746343; ROM4[526]<=26'd23452461;
ROM1[527]<=26'd1940500; ROM2[527]<=26'd11276820; ROM3[527]<=26'd9746303; ROM4[527]<=26'd23449813;
ROM1[528]<=26'd1946509; ROM2[528]<=26'd11287754; ROM3[528]<=26'd9760958; ROM4[528]<=26'd23462951;
ROM1[529]<=26'd1939975; ROM2[529]<=26'd11285435; ROM3[529]<=26'd9762602; ROM4[529]<=26'd23461337;
ROM1[530]<=26'd1929334; ROM2[530]<=26'd11280031; ROM3[530]<=26'd9759343; ROM4[530]<=26'd23455107;
ROM1[531]<=26'd1932013; ROM2[531]<=26'd11282075; ROM3[531]<=26'd9759304; ROM4[531]<=26'd23456227;
ROM1[532]<=26'd1939271; ROM2[532]<=26'd11283835; ROM3[532]<=26'd9752950; ROM4[532]<=26'd23454396;
ROM1[533]<=26'd1954776; ROM2[533]<=26'd11288931; ROM3[533]<=26'd9748862; ROM4[533]<=26'd23456442;
ROM1[534]<=26'd1959189; ROM2[534]<=26'd11290423; ROM3[534]<=26'd9749580; ROM4[534]<=26'd23459125;
ROM1[535]<=26'd1950166; ROM2[535]<=26'd11286550; ROM3[535]<=26'd9748924; ROM4[535]<=26'd23456853;
ROM1[536]<=26'd1938009; ROM2[536]<=26'd11279048; ROM3[536]<=26'd9746991; ROM4[536]<=26'd23450609;
ROM1[537]<=26'd1928073; ROM2[537]<=26'd11274123; ROM3[537]<=26'd9745652; ROM4[537]<=26'd23444636;
ROM1[538]<=26'd1922871; ROM2[538]<=26'd11276431; ROM3[538]<=26'd9748527; ROM4[538]<=26'd23446019;
ROM1[539]<=26'd1921673; ROM2[539]<=26'd11278988; ROM3[539]<=26'd9749879; ROM4[539]<=26'd23447565;
ROM1[540]<=26'd1929321; ROM2[540]<=26'd11280563; ROM3[540]<=26'd9746289; ROM4[540]<=26'd23449063;
ROM1[541]<=26'd1945464; ROM2[541]<=26'd11284827; ROM3[541]<=26'd9740534; ROM4[541]<=26'd23451371;
ROM1[542]<=26'd1953506; ROM2[542]<=26'd11285404; ROM3[542]<=26'd9736635; ROM4[542]<=26'd23450503;
ROM1[543]<=26'd1947450; ROM2[543]<=26'd11282297; ROM3[543]<=26'd9736543; ROM4[543]<=26'd23448336;
ROM1[544]<=26'd1939560; ROM2[544]<=26'd11281524; ROM3[544]<=26'd9739531; ROM4[544]<=26'd23447504;
ROM1[545]<=26'd1930546; ROM2[545]<=26'd11278608; ROM3[545]<=26'd9742539; ROM4[545]<=26'd23445899;
ROM1[546]<=26'd1925870; ROM2[546]<=26'd11279991; ROM3[546]<=26'd9748421; ROM4[546]<=26'd23449684;
ROM1[547]<=26'd1926346; ROM2[547]<=26'd11282412; ROM3[547]<=26'd9753927; ROM4[547]<=26'd23454198;
ROM1[548]<=26'd1930020; ROM2[548]<=26'd11280773; ROM3[548]<=26'd9753653; ROM4[548]<=26'd23452615;
ROM1[549]<=26'd1941399; ROM2[549]<=26'd11281252; ROM3[549]<=26'd9749707; ROM4[549]<=26'd23451913;
ROM1[550]<=26'd1951722; ROM2[550]<=26'd11282865; ROM3[550]<=26'd9746855; ROM4[550]<=26'd23452430;
ROM1[551]<=26'd1951072; ROM2[551]<=26'd11284021; ROM3[551]<=26'd9748787; ROM4[551]<=26'd23452833;
ROM1[552]<=26'd1944327; ROM2[552]<=26'd11285539; ROM3[552]<=26'd9751282; ROM4[552]<=26'd23454736;
ROM1[553]<=26'd1932097; ROM2[553]<=26'd11280928; ROM3[553]<=26'd9751844; ROM4[553]<=26'd23451324;
ROM1[554]<=26'd1924508; ROM2[554]<=26'd11279048; ROM3[554]<=26'd9754261; ROM4[554]<=26'd23448771;
ROM1[555]<=26'd1920533; ROM2[555]<=26'd11277896; ROM3[555]<=26'd9756239; ROM4[555]<=26'd23447909;
ROM1[556]<=26'd1924955; ROM2[556]<=26'd11278741; ROM3[556]<=26'd9756223; ROM4[556]<=26'd23447663;
ROM1[557]<=26'd1938454; ROM2[557]<=26'd11281601; ROM3[557]<=26'd9754718; ROM4[557]<=26'd23450373;
ROM1[558]<=26'd1949293; ROM2[558]<=26'd11279778; ROM3[558]<=26'd9749046; ROM4[558]<=26'd23449723;
ROM1[559]<=26'd1948306; ROM2[559]<=26'd11279401; ROM3[559]<=26'd9746869; ROM4[559]<=26'd23448764;
ROM1[560]<=26'd1942725; ROM2[560]<=26'd11279702; ROM3[560]<=26'd9751007; ROM4[560]<=26'd23449984;
ROM1[561]<=26'd1936457; ROM2[561]<=26'd11279223; ROM3[561]<=26'd9753759; ROM4[561]<=26'd23448867;
ROM1[562]<=26'd1930815; ROM2[562]<=26'd11278130; ROM3[562]<=26'd9752782; ROM4[562]<=26'd23445987;
ROM1[563]<=26'd1924109; ROM2[563]<=26'd11276338; ROM3[563]<=26'd9752803; ROM4[563]<=26'd23445328;
ROM1[564]<=26'd1924532; ROM2[564]<=26'd11279265; ROM3[564]<=26'd9755418; ROM4[564]<=26'd23447322;
ROM1[565]<=26'd1931785; ROM2[565]<=26'd11282321; ROM3[565]<=26'd9754686; ROM4[565]<=26'd23449568;
ROM1[566]<=26'd1944120; ROM2[566]<=26'd11281404; ROM3[566]<=26'd9748859; ROM4[566]<=26'd23448872;
ROM1[567]<=26'd1952714; ROM2[567]<=26'd11285226; ROM3[567]<=26'd9749112; ROM4[567]<=26'd23451306;
ROM1[568]<=26'd1950044; ROM2[568]<=26'd11286275; ROM3[568]<=26'd9751133; ROM4[568]<=26'd23452931;
ROM1[569]<=26'd1944876; ROM2[569]<=26'd11284241; ROM3[569]<=26'd9754848; ROM4[569]<=26'd23454971;
ROM1[570]<=26'd1936940; ROM2[570]<=26'd11282237; ROM3[570]<=26'd9757739; ROM4[570]<=26'd23455130;
ROM1[571]<=26'd1930060; ROM2[571]<=26'd11279996; ROM3[571]<=26'd9760082; ROM4[571]<=26'd23455138;
ROM1[572]<=26'd1924648; ROM2[572]<=26'd11278285; ROM3[572]<=26'd9759520; ROM4[572]<=26'd23454166;
ROM1[573]<=26'd1929847; ROM2[573]<=26'd11282165; ROM3[573]<=26'd9760102; ROM4[573]<=26'd23454233;
ROM1[574]<=26'd1948015; ROM2[574]<=26'd11288174; ROM3[574]<=26'd9761375; ROM4[574]<=26'd23458413;
ROM1[575]<=26'd1960097; ROM2[575]<=26'd11287441; ROM3[575]<=26'd9757783; ROM4[575]<=26'd23459365;
ROM1[576]<=26'd1960968; ROM2[576]<=26'd11288686; ROM3[576]<=26'd9760131; ROM4[576]<=26'd23461152;
ROM1[577]<=26'd1954539; ROM2[577]<=26'd11289469; ROM3[577]<=26'd9762915; ROM4[577]<=26'd23462969;
ROM1[578]<=26'd1952270; ROM2[578]<=26'd11295076; ROM3[578]<=26'd9771735; ROM4[578]<=26'd23469083;
ROM1[579]<=26'd1952011; ROM2[579]<=26'd11300822; ROM3[579]<=26'd9779003; ROM4[579]<=26'd23474016;
ROM1[580]<=26'd1940517; ROM2[580]<=26'd11291350; ROM3[580]<=26'd9772168; ROM4[580]<=26'd23466899;
ROM1[581]<=26'd1930840; ROM2[581]<=26'd11279145; ROM3[581]<=26'd9760394; ROM4[581]<=26'd23455410;
ROM1[582]<=26'd1936389; ROM2[582]<=26'd11275190; ROM3[582]<=26'd9753695; ROM4[582]<=26'd23451490;
ROM1[583]<=26'd1947760; ROM2[583]<=26'd11275919; ROM3[583]<=26'd9747134; ROM4[583]<=26'd23450708;
ROM1[584]<=26'd1954841; ROM2[584]<=26'd11281162; ROM3[584]<=26'd9749194; ROM4[584]<=26'd23453434;
ROM1[585]<=26'd1958010; ROM2[585]<=26'd11288464; ROM3[585]<=26'd9758020; ROM4[585]<=26'd23460191;
ROM1[586]<=26'd1953902; ROM2[586]<=26'd11292502; ROM3[586]<=26'd9763335; ROM4[586]<=26'd23462525;
ROM1[587]<=26'd1945862; ROM2[587]<=26'd11289849; ROM3[587]<=26'd9763285; ROM4[587]<=26'd23458791;
ROM1[588]<=26'd1934522; ROM2[588]<=26'd11284663; ROM3[588]<=26'd9760315; ROM4[588]<=26'd23455230;
ROM1[589]<=26'd1932742; ROM2[589]<=26'd11283066; ROM3[589]<=26'd9759015; ROM4[589]<=26'd23454131;
ROM1[590]<=26'd1933615; ROM2[590]<=26'd11279030; ROM3[590]<=26'd9749942; ROM4[590]<=26'd23448225;
ROM1[591]<=26'd1944412; ROM2[591]<=26'd11279435; ROM3[591]<=26'd9743377; ROM4[591]<=26'd23446952;
ROM1[592]<=26'd1950467; ROM2[592]<=26'd11281360; ROM3[592]<=26'd9741817; ROM4[592]<=26'd23448769;
ROM1[593]<=26'd1945992; ROM2[593]<=26'd11281616; ROM3[593]<=26'd9742747; ROM4[593]<=26'd23448837;
ROM1[594]<=26'd1941675; ROM2[594]<=26'd11283929; ROM3[594]<=26'd9746924; ROM4[594]<=26'd23452486;
ROM1[595]<=26'd1937771; ROM2[595]<=26'd11285538; ROM3[595]<=26'd9751505; ROM4[595]<=26'd23455240;
ROM1[596]<=26'd1933062; ROM2[596]<=26'd11286388; ROM3[596]<=26'd9755624; ROM4[596]<=26'd23454990;
ROM1[597]<=26'd1928480; ROM2[597]<=26'd11285994; ROM3[597]<=26'd9755275; ROM4[597]<=26'd23453449;
ROM1[598]<=26'd1932623; ROM2[598]<=26'd11285402; ROM3[598]<=26'd9752448; ROM4[598]<=26'd23452949;
ROM1[599]<=26'd1941963; ROM2[599]<=26'd11284347; ROM3[599]<=26'd9745575; ROM4[599]<=26'd23450891;
ROM1[600]<=26'd1952649; ROM2[600]<=26'd11284231; ROM3[600]<=26'd9741641; ROM4[600]<=26'd23450468;
ROM1[601]<=26'd1949470; ROM2[601]<=26'd11283074; ROM3[601]<=26'd9741147; ROM4[601]<=26'd23449717;
ROM1[602]<=26'd1938647; ROM2[602]<=26'd11278980; ROM3[602]<=26'd9740000; ROM4[602]<=26'd23444245;
ROM1[603]<=26'd1932696; ROM2[603]<=26'd11279197; ROM3[603]<=26'd9744459; ROM4[603]<=26'd23443805;
ROM1[604]<=26'd1929683; ROM2[604]<=26'd11281533; ROM3[604]<=26'd9748106; ROM4[604]<=26'd23446443;
ROM1[605]<=26'd1926035; ROM2[605]<=26'd11279929; ROM3[605]<=26'd9749919; ROM4[605]<=26'd23447023;
ROM1[606]<=26'd1930619; ROM2[606]<=26'd11283150; ROM3[606]<=26'd9752374; ROM4[606]<=26'd23448997;
ROM1[607]<=26'd1944083; ROM2[607]<=26'd11288442; ROM3[607]<=26'd9750313; ROM4[607]<=26'd23452054;
ROM1[608]<=26'd1960448; ROM2[608]<=26'd11292540; ROM3[608]<=26'd9748184; ROM4[608]<=26'd23455235;
ROM1[609]<=26'd1964513; ROM2[609]<=26'd11293879; ROM3[609]<=26'd9748102; ROM4[609]<=26'd23456112;
ROM1[610]<=26'd1950276; ROM2[610]<=26'd11285770; ROM3[610]<=26'd9741653; ROM4[610]<=26'd23449862;
ROM1[611]<=26'd1937146; ROM2[611]<=26'd11279566; ROM3[611]<=26'd9741161; ROM4[611]<=26'd23445464;
ROM1[612]<=26'd1930262; ROM2[612]<=26'd11278220; ROM3[612]<=26'd9742464; ROM4[612]<=26'd23445027;
ROM1[613]<=26'd1924771; ROM2[613]<=26'd11280577; ROM3[613]<=26'd9746063; ROM4[613]<=26'd23447451;
ROM1[614]<=26'd1929102; ROM2[614]<=26'd11284039; ROM3[614]<=26'd9751609; ROM4[614]<=26'd23452578;
ROM1[615]<=26'd1938994; ROM2[615]<=26'd11283534; ROM3[615]<=26'd9747871; ROM4[615]<=26'd23452416;
ROM1[616]<=26'd1950042; ROM2[616]<=26'd11281751; ROM3[616]<=26'd9739851; ROM4[616]<=26'd23450119;
ROM1[617]<=26'd1959462; ROM2[617]<=26'd11286590; ROM3[617]<=26'd9740966; ROM4[617]<=26'd23453441;
ROM1[618]<=26'd1957417; ROM2[618]<=26'd11291345; ROM3[618]<=26'd9746597; ROM4[618]<=26'd23456666;
ROM1[619]<=26'd1950066; ROM2[619]<=26'd11292051; ROM3[619]<=26'd9752004; ROM4[619]<=26'd23458682;
ROM1[620]<=26'd1949295; ROM2[620]<=26'd11295564; ROM3[620]<=26'd9760729; ROM4[620]<=26'd23462674;
ROM1[621]<=26'd1937168; ROM2[621]<=26'd11287424; ROM3[621]<=26'd9759083; ROM4[621]<=26'd23457070;
ROM1[622]<=26'd1925936; ROM2[622]<=26'd11278484; ROM3[622]<=26'd9753463; ROM4[622]<=26'd23451478;
ROM1[623]<=26'd1930863; ROM2[623]<=26'd11279217; ROM3[623]<=26'd9752110; ROM4[623]<=26'd23451324;
ROM1[624]<=26'd1941748; ROM2[624]<=26'd11279600; ROM3[624]<=26'd9747365; ROM4[624]<=26'd23450159;
ROM1[625]<=26'd1954637; ROM2[625]<=26'd11282612; ROM3[625]<=26'd9744223; ROM4[625]<=26'd23452872;
ROM1[626]<=26'd1958464; ROM2[626]<=26'd11286870; ROM3[626]<=26'd9748227; ROM4[626]<=26'd23457436;
ROM1[627]<=26'd1945673; ROM2[627]<=26'd11282045; ROM3[627]<=26'd9746918; ROM4[627]<=26'd23452846;
ROM1[628]<=26'd1932859; ROM2[628]<=26'd11277152; ROM3[628]<=26'd9746663; ROM4[628]<=26'd23449494;
ROM1[629]<=26'd1930186; ROM2[629]<=26'd11277250; ROM3[629]<=26'd9751364; ROM4[629]<=26'd23451917;
ROM1[630]<=26'd1927981; ROM2[630]<=26'd11278216; ROM3[630]<=26'd9753697; ROM4[630]<=26'd23451638;
ROM1[631]<=26'd1935229; ROM2[631]<=26'd11284493; ROM3[631]<=26'd9758854; ROM4[631]<=26'd23457272;
ROM1[632]<=26'd1950369; ROM2[632]<=26'd11290192; ROM3[632]<=26'd9760563; ROM4[632]<=26'd23462368;
ROM1[633]<=26'd1961486; ROM2[633]<=26'd11291270; ROM3[633]<=26'd9753619; ROM4[633]<=26'd23461680;
ROM1[634]<=26'd1963309; ROM2[634]<=26'd11292851; ROM3[634]<=26'd9751768; ROM4[634]<=26'd23463686;
ROM1[635]<=26'd1956043; ROM2[635]<=26'd11291854; ROM3[635]<=26'd9752593; ROM4[635]<=26'd23463480;
ROM1[636]<=26'd1941619; ROM2[636]<=26'd11286023; ROM3[636]<=26'd9750998; ROM4[636]<=26'd23457176;
ROM1[637]<=26'd1932459; ROM2[637]<=26'd11282472; ROM3[637]<=26'd9751713; ROM4[637]<=26'd23453619;
ROM1[638]<=26'd1928082; ROM2[638]<=26'd11281578; ROM3[638]<=26'd9756038; ROM4[638]<=26'd23454056;
ROM1[639]<=26'd1929897; ROM2[639]<=26'd11281736; ROM3[639]<=26'd9757155; ROM4[639]<=26'd23455832;
ROM1[640]<=26'd1939261; ROM2[640]<=26'd11285529; ROM3[640]<=26'd9756256; ROM4[640]<=26'd23459053;
ROM1[641]<=26'd1958117; ROM2[641]<=26'd11295028; ROM3[641]<=26'd9755968; ROM4[641]<=26'd23465877;
ROM1[642]<=26'd1964278; ROM2[642]<=26'd11296788; ROM3[642]<=26'd9751432; ROM4[642]<=26'd23464537;
ROM1[643]<=26'd1953189; ROM2[643]<=26'd11289703; ROM3[643]<=26'd9743665; ROM4[643]<=26'd23455227;
ROM1[644]<=26'd1945396; ROM2[644]<=26'd11286961; ROM3[644]<=26'd9742767; ROM4[644]<=26'd23452687;
ROM1[645]<=26'd1938866; ROM2[645]<=26'd11283973; ROM3[645]<=26'd9745334; ROM4[645]<=26'd23452880;
ROM1[646]<=26'd1932975; ROM2[646]<=26'd11283577; ROM3[646]<=26'd9749455; ROM4[646]<=26'd23454025;
ROM1[647]<=26'd1931958; ROM2[647]<=26'd11285287; ROM3[647]<=26'd9752646; ROM4[647]<=26'd23456041;
ROM1[648]<=26'd1932351; ROM2[648]<=26'd11283137; ROM3[648]<=26'd9746326; ROM4[648]<=26'd23453063;
ROM1[649]<=26'd1941942; ROM2[649]<=26'd11283839; ROM3[649]<=26'd9739071; ROM4[649]<=26'd23449416;
ROM1[650]<=26'd1952719; ROM2[650]<=26'd11284206; ROM3[650]<=26'd9736768; ROM4[650]<=26'd23449299;
ROM1[651]<=26'd1951327; ROM2[651]<=26'd11283512; ROM3[651]<=26'd9737028; ROM4[651]<=26'd23450517;
ROM1[652]<=26'd1949445; ROM2[652]<=26'd11286476; ROM3[652]<=26'd9744631; ROM4[652]<=26'd23455384;
ROM1[653]<=26'd1940824; ROM2[653]<=26'd11283259; ROM3[653]<=26'd9748380; ROM4[653]<=26'd23453432;
ROM1[654]<=26'd1933732; ROM2[654]<=26'd11278977; ROM3[654]<=26'd9747340; ROM4[654]<=26'd23450685;
ROM1[655]<=26'd1936401; ROM2[655]<=26'd11283440; ROM3[655]<=26'd9756756; ROM4[655]<=26'd23456525;
ROM1[656]<=26'd1942057; ROM2[656]<=26'd11288209; ROM3[656]<=26'd9760885; ROM4[656]<=26'd23459747;
ROM1[657]<=26'd1950842; ROM2[657]<=26'd11288007; ROM3[657]<=26'd9754024; ROM4[657]<=26'd23457536;
ROM1[658]<=26'd1961741; ROM2[658]<=26'd11287785; ROM3[658]<=26'd9746869; ROM4[658]<=26'd23455040;
ROM1[659]<=26'd1963057; ROM2[659]<=26'd11288713; ROM3[659]<=26'd9747146; ROM4[659]<=26'd23455846;
ROM1[660]<=26'd1951391; ROM2[660]<=26'd11283084; ROM3[660]<=26'd9746458; ROM4[660]<=26'd23452285;
ROM1[661]<=26'd1940938; ROM2[661]<=26'd11279707; ROM3[661]<=26'd9747469; ROM4[661]<=26'd23450920;
ROM1[662]<=26'd1940214; ROM2[662]<=26'd11284398; ROM3[662]<=26'd9755196; ROM4[662]<=26'd23456993;
ROM1[663]<=26'd1936927; ROM2[663]<=26'd11284983; ROM3[663]<=26'd9758554; ROM4[663]<=26'd23457128;
ROM1[664]<=26'd1934057; ROM2[664]<=26'd11282324; ROM3[664]<=26'd9752919; ROM4[664]<=26'd23452484;
ROM1[665]<=26'd1937941; ROM2[665]<=26'd11280654; ROM3[665]<=26'd9745835; ROM4[665]<=26'd23449969;
ROM1[666]<=26'd1947855; ROM2[666]<=26'd11280173; ROM3[666]<=26'd9736682; ROM4[666]<=26'd23444933;
ROM1[667]<=26'd1950133; ROM2[667]<=26'd11278320; ROM3[667]<=26'd9729135; ROM4[667]<=26'd23441925;
ROM1[668]<=26'd1945065; ROM2[668]<=26'd11278256; ROM3[668]<=26'd9732864; ROM4[668]<=26'd23443884;
ROM1[669]<=26'd1939248; ROM2[669]<=26'd11280679; ROM3[669]<=26'd9739753; ROM4[669]<=26'd23447373;
ROM1[670]<=26'd1934704; ROM2[670]<=26'd11280048; ROM3[670]<=26'd9744590; ROM4[670]<=26'd23450483;
ROM1[671]<=26'd1928136; ROM2[671]<=26'd11276987; ROM3[671]<=26'd9745481; ROM4[671]<=26'd23448008;
ROM1[672]<=26'd1927076; ROM2[672]<=26'd11279134; ROM3[672]<=26'd9745750; ROM4[672]<=26'd23448507;
ROM1[673]<=26'd1935546; ROM2[673]<=26'd11282024; ROM3[673]<=26'd9746032; ROM4[673]<=26'd23449520;
ROM1[674]<=26'd1940605; ROM2[674]<=26'd11278302; ROM3[674]<=26'd9738217; ROM4[674]<=26'd23442961;
ROM1[675]<=26'd1945367; ROM2[675]<=26'd11276725; ROM3[675]<=26'd9732414; ROM4[675]<=26'd23440666;
ROM1[676]<=26'd1946036; ROM2[676]<=26'd11276407; ROM3[676]<=26'd9734607; ROM4[676]<=26'd23441782;
ROM1[677]<=26'd1938848; ROM2[677]<=26'd11273952; ROM3[677]<=26'd9735765; ROM4[677]<=26'd23440162;
ROM1[678]<=26'd1929625; ROM2[678]<=26'd11270555; ROM3[678]<=26'd9735087; ROM4[678]<=26'd23437332;
ROM1[679]<=26'd1920873; ROM2[679]<=26'd11269575; ROM3[679]<=26'd9735976; ROM4[679]<=26'd23435712;
ROM1[680]<=26'd1915235; ROM2[680]<=26'd11268701; ROM3[680]<=26'd9738087; ROM4[680]<=26'd23434473;
ROM1[681]<=26'd1917108; ROM2[681]<=26'd11268683; ROM3[681]<=26'd9737812; ROM4[681]<=26'd23432669;
ROM1[682]<=26'd1931575; ROM2[682]<=26'd11274144; ROM3[682]<=26'd9738339; ROM4[682]<=26'd23437070;
ROM1[683]<=26'd1950957; ROM2[683]<=26'd11280986; ROM3[683]<=26'd9737328; ROM4[683]<=26'd23443296;
ROM1[684]<=26'd1954534; ROM2[684]<=26'd11282363; ROM3[684]<=26'd9739452; ROM4[684]<=26'd23446093;
ROM1[685]<=26'd1946468; ROM2[685]<=26'd11280209; ROM3[685]<=26'd9741320; ROM4[685]<=26'd23446621;
ROM1[686]<=26'd1947747; ROM2[686]<=26'd11289174; ROM3[686]<=26'd9754190; ROM4[686]<=26'd23457226;
ROM1[687]<=26'd1952451; ROM2[687]<=26'd11296236; ROM3[687]<=26'd9767289; ROM4[687]<=26'd23466584;
ROM1[688]<=26'd1936184; ROM2[688]<=26'd11284857; ROM3[688]<=26'd9757163; ROM4[688]<=26'd23455979;
ROM1[689]<=26'd1926619; ROM2[689]<=26'd11275008; ROM3[689]<=26'd9748221; ROM4[689]<=26'd23447795;
ROM1[690]<=26'd1932472; ROM2[690]<=26'd11274405; ROM3[690]<=26'd9744990; ROM4[690]<=26'd23446901;
ROM1[691]<=26'd1940717; ROM2[691]<=26'd11273603; ROM3[691]<=26'd9737961; ROM4[691]<=26'd23443896;
ROM1[692]<=26'd1949857; ROM2[692]<=26'd11275986; ROM3[692]<=26'd9740227; ROM4[692]<=26'd23447549;
ROM1[693]<=26'd1952524; ROM2[693]<=26'd11282011; ROM3[693]<=26'd9749129; ROM4[693]<=26'd23456246;
ROM1[694]<=26'd1945047; ROM2[694]<=26'd11281492; ROM3[694]<=26'd9753566; ROM4[694]<=26'd23457703;
ROM1[695]<=26'd1942057; ROM2[695]<=26'd11284554; ROM3[695]<=26'd9758330; ROM4[695]<=26'd23460273;
ROM1[696]<=26'd1941324; ROM2[696]<=26'd11289847; ROM3[696]<=26'd9764565; ROM4[696]<=26'd23466897;
ROM1[697]<=26'd1939471; ROM2[697]<=26'd11290501; ROM3[697]<=26'd9766692; ROM4[697]<=26'd23467597;
ROM1[698]<=26'd1942795; ROM2[698]<=26'd11290430; ROM3[698]<=26'd9764363; ROM4[698]<=26'd23466773;
ROM1[699]<=26'd1952145; ROM2[699]<=26'd11287791; ROM3[699]<=26'd9757226; ROM4[699]<=26'd23463553;
ROM1[700]<=26'd1970221; ROM2[700]<=26'd11296675; ROM3[700]<=26'd9760475; ROM4[700]<=26'd23469752;
ROM1[701]<=26'd1971799; ROM2[701]<=26'd11300748; ROM3[701]<=26'd9761844; ROM4[701]<=26'd23473059;
ROM1[702]<=26'd1957813; ROM2[702]<=26'd11293194; ROM3[702]<=26'd9754663; ROM4[702]<=26'd23464545;
ROM1[703]<=26'd1948211; ROM2[703]<=26'd11289373; ROM3[703]<=26'd9753106; ROM4[703]<=26'd23459865;
ROM1[704]<=26'd1943178; ROM2[704]<=26'd11289045; ROM3[704]<=26'd9755392; ROM4[704]<=26'd23459719;
ROM1[705]<=26'd1937986; ROM2[705]<=26'd11288891; ROM3[705]<=26'd9759012; ROM4[705]<=26'd23458690;
ROM1[706]<=26'd1938918; ROM2[706]<=26'd11286833; ROM3[706]<=26'd9756336; ROM4[706]<=26'd23456064;
ROM1[707]<=26'd1948534; ROM2[707]<=26'd11288757; ROM3[707]<=26'd9751349; ROM4[707]<=26'd23457980;
ROM1[708]<=26'd1959787; ROM2[708]<=26'd11290436; ROM3[708]<=26'd9745397; ROM4[708]<=26'd23457328;
ROM1[709]<=26'd1964064; ROM2[709]<=26'd11292488; ROM3[709]<=26'd9745614; ROM4[709]<=26'd23458366;
ROM1[710]<=26'd1962420; ROM2[710]<=26'd11296357; ROM3[710]<=26'd9752187; ROM4[710]<=26'd23463592;
ROM1[711]<=26'd1957900; ROM2[711]<=26'd11297649; ROM3[711]<=26'd9757232; ROM4[711]<=26'd23467087;
ROM1[712]<=26'd1951112; ROM2[712]<=26'd11295517; ROM3[712]<=26'd9757925; ROM4[712]<=26'd23466209;
ROM1[713]<=26'd1942216; ROM2[713]<=26'd11291610; ROM3[713]<=26'd9757857; ROM4[713]<=26'd23462538;
ROM1[714]<=26'd1940480; ROM2[714]<=26'd11290477; ROM3[714]<=26'd9756622; ROM4[714]<=26'd23461673;
ROM1[715]<=26'd1943516; ROM2[715]<=26'd11289032; ROM3[715]<=26'd9751364; ROM4[715]<=26'd23458048;
ROM1[716]<=26'd1952844; ROM2[716]<=26'd11286578; ROM3[716]<=26'd9741688; ROM4[716]<=26'd23454400;
ROM1[717]<=26'd1957362; ROM2[717]<=26'd11285112; ROM3[717]<=26'd9735756; ROM4[717]<=26'd23452850;
ROM1[718]<=26'd1952159; ROM2[718]<=26'd11284774; ROM3[718]<=26'd9735458; ROM4[718]<=26'd23451659;
ROM1[719]<=26'd1944659; ROM2[719]<=26'd11283492; ROM3[719]<=26'd9735885; ROM4[719]<=26'd23448794;
ROM1[720]<=26'd1936737; ROM2[720]<=26'd11282457; ROM3[720]<=26'd9737000; ROM4[720]<=26'd23445800;
ROM1[721]<=26'd1928561; ROM2[721]<=26'd11282347; ROM3[721]<=26'd9741027; ROM4[721]<=26'd23445232;
ROM1[722]<=26'd1924896; ROM2[722]<=26'd11281019; ROM3[722]<=26'd9742521; ROM4[722]<=26'd23445330;
ROM1[723]<=26'd1929062; ROM2[723]<=26'd11280558; ROM3[723]<=26'd9741436; ROM4[723]<=26'd23445598;
ROM1[724]<=26'd1941859; ROM2[724]<=26'd11283137; ROM3[724]<=26'd9739350; ROM4[724]<=26'd23446493;
ROM1[725]<=26'd1956710; ROM2[725]<=26'd11288225; ROM3[725]<=26'd9737193; ROM4[725]<=26'd23450597;
ROM1[726]<=26'd1957457; ROM2[726]<=26'd11290644; ROM3[726]<=26'd9738189; ROM4[726]<=26'd23452264;
ROM1[727]<=26'd1948322; ROM2[727]<=26'd11286761; ROM3[727]<=26'd9739535; ROM4[727]<=26'd23450672;
ROM1[728]<=26'd1939959; ROM2[728]<=26'd11284818; ROM3[728]<=26'd9743806; ROM4[728]<=26'd23450064;
ROM1[729]<=26'd1937333; ROM2[729]<=26'd11287686; ROM3[729]<=26'd9751836; ROM4[729]<=26'd23454827;
ROM1[730]<=26'd1935761; ROM2[730]<=26'd11290727; ROM3[730]<=26'd9760285; ROM4[730]<=26'd23459262;
ROM1[731]<=26'd1936742; ROM2[731]<=26'd11291253; ROM3[731]<=26'd9757541; ROM4[731]<=26'd23457064;
ROM1[732]<=26'd1944555; ROM2[732]<=26'd11289376; ROM3[732]<=26'd9750342; ROM4[732]<=26'd23452835;
ROM1[733]<=26'd1952679; ROM2[733]<=26'd11286644; ROM3[733]<=26'd9741967; ROM4[733]<=26'd23449293;
ROM1[734]<=26'd1952991; ROM2[734]<=26'd11284063; ROM3[734]<=26'd9740345; ROM4[734]<=26'd23449103;
ROM1[735]<=26'd1951804; ROM2[735]<=26'd11286984; ROM3[735]<=26'd9749319; ROM4[735]<=26'd23454359;
ROM1[736]<=26'd1955084; ROM2[736]<=26'd11298367; ROM3[736]<=26'd9763640; ROM4[736]<=26'd23465664;
ROM1[737]<=26'd1960899; ROM2[737]<=26'd11307400; ROM3[737]<=26'd9775123; ROM4[737]<=26'd23474319;
ROM1[738]<=26'd1952514; ROM2[738]<=26'd11302082; ROM3[738]<=26'd9772591; ROM4[738]<=26'd23469629;
ROM1[739]<=26'd1941029; ROM2[739]<=26'd11291512; ROM3[739]<=26'd9764485; ROM4[739]<=26'd23459865;
ROM1[740]<=26'd1941165; ROM2[740]<=26'd11284501; ROM3[740]<=26'd9755229; ROM4[740]<=26'd23452976;
ROM1[741]<=26'd1951759; ROM2[741]<=26'd11284173; ROM3[741]<=26'd9748485; ROM4[741]<=26'd23452190;
ROM1[742]<=26'd1966069; ROM2[742]<=26'd11294160; ROM3[742]<=26'd9753561; ROM4[742]<=26'd23460258;
ROM1[743]<=26'd1968161; ROM2[743]<=26'd11299754; ROM3[743]<=26'd9761337; ROM4[743]<=26'd23465944;
ROM1[744]<=26'd1954210; ROM2[744]<=26'd11291758; ROM3[744]<=26'd9759936; ROM4[744]<=26'd23461198;
ROM1[745]<=26'd1945809; ROM2[745]<=26'd11288446; ROM3[745]<=26'd9760727; ROM4[745]<=26'd23459333;
ROM1[746]<=26'd1938044; ROM2[746]<=26'd11285269; ROM3[746]<=26'd9761951; ROM4[746]<=26'd23459615;
ROM1[747]<=26'd1937620; ROM2[747]<=26'd11287540; ROM3[747]<=26'd9763465; ROM4[747]<=26'd23463187;
ROM1[748]<=26'd1953036; ROM2[748]<=26'd11299089; ROM3[748]<=26'd9770222; ROM4[748]<=26'd23471813;
ROM1[749]<=26'd1962840; ROM2[749]<=26'd11297217; ROM3[749]<=26'd9763709; ROM4[749]<=26'd23468002;
ROM1[750]<=26'd1968922; ROM2[750]<=26'd11294172; ROM3[750]<=26'd9756053; ROM4[750]<=26'd23463192;
ROM1[751]<=26'd1972743; ROM2[751]<=26'd11300427; ROM3[751]<=26'd9762810; ROM4[751]<=26'd23470437;
ROM1[752]<=26'd1964289; ROM2[752]<=26'd11296493; ROM3[752]<=26'd9764194; ROM4[752]<=26'd23470614;
ROM1[753]<=26'd1956606; ROM2[753]<=26'd11292655; ROM3[753]<=26'd9764505; ROM4[753]<=26'd23467901;
ROM1[754]<=26'd1952691; ROM2[754]<=26'd11292428; ROM3[754]<=26'd9767595; ROM4[754]<=26'd23468133;
ROM1[755]<=26'd1945375; ROM2[755]<=26'd11288048; ROM3[755]<=26'd9766271; ROM4[755]<=26'd23464505;
ROM1[756]<=26'd1947320; ROM2[756]<=26'd11288463; ROM3[756]<=26'd9764329; ROM4[756]<=26'd23465003;
ROM1[757]<=26'd1958231; ROM2[757]<=26'd11291818; ROM3[757]<=26'd9763352; ROM4[757]<=26'd23467589;
ROM1[758]<=26'd1971546; ROM2[758]<=26'd11295338; ROM3[758]<=26'd9761427; ROM4[758]<=26'd23469425;
ROM1[759]<=26'd1974139; ROM2[759]<=26'd11297344; ROM3[759]<=26'd9762754; ROM4[759]<=26'd23471174;
ROM1[760]<=26'd1964878; ROM2[760]<=26'd11293595; ROM3[760]<=26'd9762388; ROM4[760]<=26'd23467309;
ROM1[761]<=26'd1955944; ROM2[761]<=26'd11292962; ROM3[761]<=26'd9763815; ROM4[761]<=26'd23466749;
ROM1[762]<=26'd1953860; ROM2[762]<=26'd11296895; ROM3[762]<=26'd9768855; ROM4[762]<=26'd23470827;
ROM1[763]<=26'd1943118; ROM2[763]<=26'd11289913; ROM3[763]<=26'd9764985; ROM4[763]<=26'd23463313;
ROM1[764]<=26'd1938837; ROM2[764]<=26'd11286745; ROM3[764]<=26'd9760081; ROM4[764]<=26'd23459447;
ROM1[765]<=26'd1944930; ROM2[765]<=26'd11287897; ROM3[765]<=26'd9754319; ROM4[765]<=26'd23457787;
ROM1[766]<=26'd1953652; ROM2[766]<=26'd11283944; ROM3[766]<=26'd9744684; ROM4[766]<=26'd23451365;
ROM1[767]<=26'd1957020; ROM2[767]<=26'd11282413; ROM3[767]<=26'd9738407; ROM4[767]<=26'd23448264;
ROM1[768]<=26'd1951647; ROM2[768]<=26'd11281187; ROM3[768]<=26'd9740713; ROM4[768]<=26'd23448234;
ROM1[769]<=26'd1947522; ROM2[769]<=26'd11281113; ROM3[769]<=26'd9747327; ROM4[769]<=26'd23450464;
ROM1[770]<=26'd1941276; ROM2[770]<=26'd11280888; ROM3[770]<=26'd9748364; ROM4[770]<=26'd23449120;
ROM1[771]<=26'd1933788; ROM2[771]<=26'd11280262; ROM3[771]<=26'd9751441; ROM4[771]<=26'd23448821;
ROM1[772]<=26'd1938188; ROM2[772]<=26'd11286139; ROM3[772]<=26'd9760257; ROM4[772]<=26'd23456086;
ROM1[773]<=26'd1951824; ROM2[773]<=26'd11296870; ROM3[773]<=26'd9768758; ROM4[773]<=26'd23465339;
ROM1[774]<=26'd1963186; ROM2[774]<=26'd11298975; ROM3[774]<=26'd9765492; ROM4[774]<=26'd23465895;
ROM1[775]<=26'd1968439; ROM2[775]<=26'd11296143; ROM3[775]<=26'd9756470; ROM4[775]<=26'd23463117;
ROM1[776]<=26'd1961346; ROM2[776]<=26'd11293190; ROM3[776]<=26'd9753072; ROM4[776]<=26'd23459624;
ROM1[777]<=26'd1946971; ROM2[777]<=26'd11284106; ROM3[777]<=26'd9749517; ROM4[777]<=26'd23453248;
ROM1[778]<=26'd1937105; ROM2[778]<=26'd11278204; ROM3[778]<=26'd9748521; ROM4[778]<=26'd23450061;
ROM1[779]<=26'd1935702; ROM2[779]<=26'd11282261; ROM3[779]<=26'd9756576; ROM4[779]<=26'd23455690;
ROM1[780]<=26'd1933550; ROM2[780]<=26'd11284675; ROM3[780]<=26'd9761460; ROM4[780]<=26'd23458992;
ROM1[781]<=26'd1933769; ROM2[781]<=26'd11282865; ROM3[781]<=26'd9757294; ROM4[781]<=26'd23455737;
ROM1[782]<=26'd1943702; ROM2[782]<=26'd11285428; ROM3[782]<=26'd9753877; ROM4[782]<=26'd23455670;
ROM1[783]<=26'd1957086; ROM2[783]<=26'd11286799; ROM3[783]<=26'd9748380; ROM4[783]<=26'd23454831;
ROM1[784]<=26'd1961490; ROM2[784]<=26'd11288042; ROM3[784]<=26'd9749622; ROM4[784]<=26'd23458077;
ROM1[785]<=26'd1956817; ROM2[785]<=26'd11289244; ROM3[785]<=26'd9754603; ROM4[785]<=26'd23460730;
ROM1[786]<=26'd1950031; ROM2[786]<=26'd11289290; ROM3[786]<=26'd9757923; ROM4[786]<=26'd23462531;
ROM1[787]<=26'd1947998; ROM2[787]<=26'd11292326; ROM3[787]<=26'd9763876; ROM4[787]<=26'd23466199;
ROM1[788]<=26'd1945748; ROM2[788]<=26'd11295280; ROM3[788]<=26'd9767399; ROM4[788]<=26'd23467377;
ROM1[789]<=26'd1942075; ROM2[789]<=26'd11291363; ROM3[789]<=26'd9761937; ROM4[789]<=26'd23461576;
ROM1[790]<=26'd1945822; ROM2[790]<=26'd11289042; ROM3[790]<=26'd9755378; ROM4[790]<=26'd23458264;
ROM1[791]<=26'd1958601; ROM2[791]<=26'd11291936; ROM3[791]<=26'd9749262; ROM4[791]<=26'd23458062;
ROM1[792]<=26'd1962692; ROM2[792]<=26'd11291256; ROM3[792]<=26'd9742108; ROM4[792]<=26'd23453640;
ROM1[793]<=26'd1956359; ROM2[793]<=26'd11292384; ROM3[793]<=26'd9742811; ROM4[793]<=26'd23454727;
ROM1[794]<=26'd1948829; ROM2[794]<=26'd11295395; ROM3[794]<=26'd9748195; ROM4[794]<=26'd23456370;
ROM1[795]<=26'd1942338; ROM2[795]<=26'd11293970; ROM3[795]<=26'd9750576; ROM4[795]<=26'd23454710;
ROM1[796]<=26'd1935127; ROM2[796]<=26'd11292687; ROM3[796]<=26'd9753495; ROM4[796]<=26'd23455427;
ROM1[797]<=26'd1934764; ROM2[797]<=26'd11293190; ROM3[797]<=26'd9756670; ROM4[797]<=26'd23456798;
ROM1[798]<=26'd1940985; ROM2[798]<=26'd11291728; ROM3[798]<=26'd9756149; ROM4[798]<=26'd23455727;
ROM1[799]<=26'd1953373; ROM2[799]<=26'd11291463; ROM3[799]<=26'd9752570; ROM4[799]<=26'd23456439;
ROM1[800]<=26'd1959446; ROM2[800]<=26'd11289335; ROM3[800]<=26'd9746222; ROM4[800]<=26'd23453530;
ROM1[801]<=26'd1952929; ROM2[801]<=26'd11284770; ROM3[801]<=26'd9742130; ROM4[801]<=26'd23448586;
ROM1[802]<=26'd1946943; ROM2[802]<=26'd11283798; ROM3[802]<=26'd9745662; ROM4[802]<=26'd23449749;
ROM1[803]<=26'd1939707; ROM2[803]<=26'd11282716; ROM3[803]<=26'd9748188; ROM4[803]<=26'd23449749;
ROM1[804]<=26'd1935481; ROM2[804]<=26'd11283749; ROM3[804]<=26'd9753003; ROM4[804]<=26'd23452783;
ROM1[805]<=26'd1932315; ROM2[805]<=26'd11284738; ROM3[805]<=26'd9757486; ROM4[805]<=26'd23455786;
ROM1[806]<=26'd1932686; ROM2[806]<=26'd11282991; ROM3[806]<=26'd9754350; ROM4[806]<=26'd23455402;
ROM1[807]<=26'd1941324; ROM2[807]<=26'd11285126; ROM3[807]<=26'd9752398; ROM4[807]<=26'd23455796;
ROM1[808]<=26'd1954034; ROM2[808]<=26'd11285981; ROM3[808]<=26'd9746355; ROM4[808]<=26'd23454567;
ROM1[809]<=26'd1956586; ROM2[809]<=26'd11287364; ROM3[809]<=26'd9745582; ROM4[809]<=26'd23455632;
ROM1[810]<=26'd1952269; ROM2[810]<=26'd11290794; ROM3[810]<=26'd9751538; ROM4[810]<=26'd23458786;
ROM1[811]<=26'd1949063; ROM2[811]<=26'd11291836; ROM3[811]<=26'd9756799; ROM4[811]<=26'd23462419;
ROM1[812]<=26'd1947182; ROM2[812]<=26'd11294870; ROM3[812]<=26'd9760423; ROM4[812]<=26'd23466880;
ROM1[813]<=26'd1944842; ROM2[813]<=26'd11296634; ROM3[813]<=26'd9765346; ROM4[813]<=26'd23470075;
ROM1[814]<=26'd1944925; ROM2[814]<=26'd11296555; ROM3[814]<=26'd9766058; ROM4[814]<=26'd23469709;
ROM1[815]<=26'd1948189; ROM2[815]<=26'd11294093; ROM3[815]<=26'd9760663; ROM4[815]<=26'd23466261;
ROM1[816]<=26'd1958223; ROM2[816]<=26'd11293114; ROM3[816]<=26'd9754694; ROM4[816]<=26'd23462818;
ROM1[817]<=26'd1957409; ROM2[817]<=26'd11289702; ROM3[817]<=26'd9745372; ROM4[817]<=26'd23458153;
ROM1[818]<=26'd1947289; ROM2[818]<=26'd11284615; ROM3[818]<=26'd9741914; ROM4[818]<=26'd23452858;
ROM1[819]<=26'd1941747; ROM2[819]<=26'd11285153; ROM3[819]<=26'd9745495; ROM4[819]<=26'd23453219;
ROM1[820]<=26'd1938774; ROM2[820]<=26'd11286283; ROM3[820]<=26'd9752338; ROM4[820]<=26'd23455570;
ROM1[821]<=26'd1934521; ROM2[821]<=26'd11286922; ROM3[821]<=26'd9759574; ROM4[821]<=26'd23458346;
ROM1[822]<=26'd1933070; ROM2[822]<=26'd11287736; ROM3[822]<=26'd9761776; ROM4[822]<=26'd23461082;
ROM1[823]<=26'd1938609; ROM2[823]<=26'd11286769; ROM3[823]<=26'd9759599; ROM4[823]<=26'd23461381;
ROM1[824]<=26'd1953582; ROM2[824]<=26'd11291381; ROM3[824]<=26'd9758981; ROM4[824]<=26'd23464760;
ROM1[825]<=26'd1960810; ROM2[825]<=26'd11292048; ROM3[825]<=26'd9755081; ROM4[825]<=26'd23463144;
ROM1[826]<=26'd1954733; ROM2[826]<=26'd11287940; ROM3[826]<=26'd9753013; ROM4[826]<=26'd23459408;
ROM1[827]<=26'd1947474; ROM2[827]<=26'd11288886; ROM3[827]<=26'd9757685; ROM4[827]<=26'd23460475;
ROM1[828]<=26'd1934454; ROM2[828]<=26'd11283830; ROM3[828]<=26'd9756640; ROM4[828]<=26'd23455603;
ROM1[829]<=26'd1926879; ROM2[829]<=26'd11281286; ROM3[829]<=26'd9756636; ROM4[829]<=26'd23452709;
ROM1[830]<=26'd1928977; ROM2[830]<=26'd11288611; ROM3[830]<=26'd9763377; ROM4[830]<=26'd23457851;
ROM1[831]<=26'd1942916; ROM2[831]<=26'd11299630; ROM3[831]<=26'd9773056; ROM4[831]<=26'd23468134;
ROM1[832]<=26'd1951760; ROM2[832]<=26'd11298256; ROM3[832]<=26'd9766073; ROM4[832]<=26'd23467107;
ROM1[833]<=26'd1957508; ROM2[833]<=26'd11292718; ROM3[833]<=26'd9754015; ROM4[833]<=26'd23460577;
ROM1[834]<=26'd1960165; ROM2[834]<=26'd11292817; ROM3[834]<=26'd9754104; ROM4[834]<=26'd23460453;
ROM1[835]<=26'd1952161; ROM2[835]<=26'd11291457; ROM3[835]<=26'd9754799; ROM4[835]<=26'd23460218;
ROM1[836]<=26'd1947377; ROM2[836]<=26'd11294973; ROM3[836]<=26'd9761598; ROM4[836]<=26'd23463630;
ROM1[837]<=26'd1944995; ROM2[837]<=26'd11297315; ROM3[837]<=26'd9764078; ROM4[837]<=26'd23465341;
ROM1[838]<=26'd1932770; ROM2[838]<=26'd11290478; ROM3[838]<=26'd9758867; ROM4[838]<=26'd23459811;
ROM1[839]<=26'd1926516; ROM2[839]<=26'd11284380; ROM3[839]<=26'd9752974; ROM4[839]<=26'd23454299;
ROM1[840]<=26'd1927873; ROM2[840]<=26'd11278117; ROM3[840]<=26'd9742736; ROM4[840]<=26'd23447921;
ROM1[841]<=26'd1940113; ROM2[841]<=26'd11280162; ROM3[841]<=26'd9737484; ROM4[841]<=26'd23447745;
ROM1[842]<=26'd1951711; ROM2[842]<=26'd11286766; ROM3[842]<=26'd9742309; ROM4[842]<=26'd23453746;
ROM1[843]<=26'd1947568; ROM2[843]<=26'd11287544; ROM3[843]<=26'd9744735; ROM4[843]<=26'd23454275;
ROM1[844]<=26'd1936794; ROM2[844]<=26'd11284695; ROM3[844]<=26'd9745206; ROM4[844]<=26'd23452044;
ROM1[845]<=26'd1929334; ROM2[845]<=26'd11281315; ROM3[845]<=26'd9747839; ROM4[845]<=26'd23450493;
ROM1[846]<=26'd1930696; ROM2[846]<=26'd11288110; ROM3[846]<=26'd9756863; ROM4[846]<=26'd23458519;
ROM1[847]<=26'd1927230; ROM2[847]<=26'd11288481; ROM3[847]<=26'd9756933; ROM4[847]<=26'd23457941;
ROM1[848]<=26'd1929719; ROM2[848]<=26'd11284922; ROM3[848]<=26'd9751682; ROM4[848]<=26'd23452878;
ROM1[849]<=26'd1943804; ROM2[849]<=26'd11287485; ROM3[849]<=26'd9748780; ROM4[849]<=26'd23455606;
ROM1[850]<=26'd1952332; ROM2[850]<=26'd11288726; ROM3[850]<=26'd9744428; ROM4[850]<=26'd23455984;
ROM1[851]<=26'd1946493; ROM2[851]<=26'd11285025; ROM3[851]<=26'd9740209; ROM4[851]<=26'd23452432;
ROM1[852]<=26'd1942095; ROM2[852]<=26'd11286629; ROM3[852]<=26'd9744792; ROM4[852]<=26'd23454038;
ROM1[853]<=26'd1943026; ROM2[853]<=26'd11290835; ROM3[853]<=26'd9755677; ROM4[853]<=26'd23460272;
ROM1[854]<=26'd1934274; ROM2[854]<=26'd11286086; ROM3[854]<=26'd9756121; ROM4[854]<=26'd23458670;
ROM1[855]<=26'd1928325; ROM2[855]<=26'd11285317; ROM3[855]<=26'd9760920; ROM4[855]<=26'd23459021;
ROM1[856]<=26'd1932317; ROM2[856]<=26'd11287336; ROM3[856]<=26'd9765997; ROM4[856]<=26'd23463068;
ROM1[857]<=26'd1944845; ROM2[857]<=26'd11291313; ROM3[857]<=26'd9765161; ROM4[857]<=26'd23466380;
ROM1[858]<=26'd1958283; ROM2[858]<=26'd11293150; ROM3[858]<=26'd9761865; ROM4[858]<=26'd23467168;
ROM1[859]<=26'd1963237; ROM2[859]<=26'd11294614; ROM3[859]<=26'd9763623; ROM4[859]<=26'd23469318;
ROM1[860]<=26'd1963748; ROM2[860]<=26'd11299634; ROM3[860]<=26'd9773638; ROM4[860]<=26'd23475383;
ROM1[861]<=26'd1954772; ROM2[861]<=26'd11298367; ROM3[861]<=26'd9777965; ROM4[861]<=26'd23475662;
ROM1[862]<=26'd1948422; ROM2[862]<=26'd11295441; ROM3[862]<=26'd9778687; ROM4[862]<=26'd23474773;
ROM1[863]<=26'd1943691; ROM2[863]<=26'd11293319; ROM3[863]<=26'd9780758; ROM4[863]<=26'd23476104;
ROM1[864]<=26'd1941021; ROM2[864]<=26'd11293188; ROM3[864]<=26'd9778079; ROM4[864]<=26'd23476254;
ROM1[865]<=26'd1957899; ROM2[865]<=26'd11303065; ROM3[865]<=26'd9781032; ROM4[865]<=26'd23485346;
ROM1[866]<=26'd1974649; ROM2[866]<=26'd11306533; ROM3[866]<=26'd9778053; ROM4[866]<=26'd23485867;
ROM1[867]<=26'd1971172; ROM2[867]<=26'd11301578; ROM3[867]<=26'd9766945; ROM4[867]<=26'd23477800;
ROM1[868]<=26'd1961085; ROM2[868]<=26'd11298860; ROM3[868]<=26'd9764715; ROM4[868]<=26'd23474472;
ROM1[869]<=26'd1957666; ROM2[869]<=26'd11297633; ROM3[869]<=26'd9767996; ROM4[869]<=26'd23474371;
ROM1[870]<=26'd1955400; ROM2[870]<=26'd11297926; ROM3[870]<=26'd9769154; ROM4[870]<=26'd23476167;
ROM1[871]<=26'd1957191; ROM2[871]<=26'd11301964; ROM3[871]<=26'd9775068; ROM4[871]<=26'd23480984;
ROM1[872]<=26'd1957810; ROM2[872]<=26'd11302951; ROM3[872]<=26'd9774200; ROM4[872]<=26'd23480421;
ROM1[873]<=26'd1958022; ROM2[873]<=26'd11301623; ROM3[873]<=26'd9768767; ROM4[873]<=26'd23477960;
ROM1[874]<=26'd1969105; ROM2[874]<=26'd11301360; ROM3[874]<=26'd9762182; ROM4[874]<=26'd23474264;
ROM1[875]<=26'd1983740; ROM2[875]<=26'd11305574; ROM3[875]<=26'd9759675; ROM4[875]<=26'd23476670;
ROM1[876]<=26'd1984820; ROM2[876]<=26'd11306001; ROM3[876]<=26'd9760988; ROM4[876]<=26'd23477962;
ROM1[877]<=26'd1969716; ROM2[877]<=26'd11296707; ROM3[877]<=26'd9754982; ROM4[877]<=26'd23467315;
ROM1[878]<=26'd1965235; ROM2[878]<=26'd11299773; ROM3[878]<=26'd9761375; ROM4[878]<=26'd23471789;
ROM1[879]<=26'd1963433; ROM2[879]<=26'd11299833; ROM3[879]<=26'd9767833; ROM4[879]<=26'd23475130;
ROM1[880]<=26'd1962484; ROM2[880]<=26'd11298013; ROM3[880]<=26'd9771745; ROM4[880]<=26'd23476679;
ROM1[881]<=26'd1972837; ROM2[881]<=26'd11304416; ROM3[881]<=26'd9777687; ROM4[881]<=26'd23483485;
ROM1[882]<=26'd1987083; ROM2[882]<=26'd11309348; ROM3[882]<=26'd9771771; ROM4[882]<=26'd23482227;
ROM1[883]<=26'd1999578; ROM2[883]<=26'd11310198; ROM3[883]<=26'd9762877; ROM4[883]<=26'd23478451;
ROM1[884]<=26'd2003438; ROM2[884]<=26'd11309301; ROM3[884]<=26'd9761005; ROM4[884]<=26'd23477853;
ROM1[885]<=26'd2003658; ROM2[885]<=26'd11313814; ROM3[885]<=26'd9767739; ROM4[885]<=26'd23482712;
ROM1[886]<=26'd2007087; ROM2[886]<=26'd11322887; ROM3[886]<=26'd9781582; ROM4[886]<=26'd23494196;
ROM1[887]<=26'd2006353; ROM2[887]<=26'd11325286; ROM3[887]<=26'd9785287; ROM4[887]<=26'd23495667;
ROM1[888]<=26'd1999874; ROM2[888]<=26'd11321355; ROM3[888]<=26'd9780727; ROM4[888]<=26'd23489131;
ROM1[889]<=26'd2011689; ROM2[889]<=26'd11327520; ROM3[889]<=26'd9785681; ROM4[889]<=26'd23493397;
ROM1[890]<=26'd2024938; ROM2[890]<=26'd11328664; ROM3[890]<=26'd9786558; ROM4[890]<=26'd23494352;
ROM1[891]<=26'd2035345; ROM2[891]<=26'd11326641; ROM3[891]<=26'd9778282; ROM4[891]<=26'd23492210;
ROM1[892]<=26'd2046739; ROM2[892]<=26'd11331991; ROM3[892]<=26'd9777897; ROM4[892]<=26'd23495905;
ROM1[893]<=26'd2045204; ROM2[893]<=26'd11331931; ROM3[893]<=26'd9776027; ROM4[893]<=26'd23495230;
ROM1[894]<=26'd2037320; ROM2[894]<=26'd11327300; ROM3[894]<=26'd9771598; ROM4[894]<=26'd23489964;
ROM1[895]<=26'd2034798; ROM2[895]<=26'd11327874; ROM3[895]<=26'd9774841; ROM4[895]<=26'd23490716;
ROM1[896]<=26'd2031407; ROM2[896]<=26'd11330796; ROM3[896]<=26'd9779880; ROM4[896]<=26'd23495120;
ROM1[897]<=26'd2029222; ROM2[897]<=26'd11329257; ROM3[897]<=26'd9779988; ROM4[897]<=26'd23494161;
ROM1[898]<=26'd2032195; ROM2[898]<=26'd11325682; ROM3[898]<=26'd9774148; ROM4[898]<=26'd23490453;
ROM1[899]<=26'd2042662; ROM2[899]<=26'd11323692; ROM3[899]<=26'd9765720; ROM4[899]<=26'd23487072;
ROM1[900]<=26'd2058239; ROM2[900]<=26'd11327150; ROM3[900]<=26'd9763752; ROM4[900]<=26'd23489887;
ROM1[901]<=26'd2056697; ROM2[901]<=26'd11328413; ROM3[901]<=26'd9763546; ROM4[901]<=26'd23491237;
ROM1[902]<=26'd2045421; ROM2[902]<=26'd11324741; ROM3[902]<=26'd9763275; ROM4[902]<=26'd23487221;
ROM1[903]<=26'd2038755; ROM2[903]<=26'd11325051; ROM3[903]<=26'd9767508; ROM4[903]<=26'd23487946;
ROM1[904]<=26'd2034030; ROM2[904]<=26'd11328233; ROM3[904]<=26'd9771884; ROM4[904]<=26'd23489312;
ROM1[905]<=26'd2028116; ROM2[905]<=26'd11326321; ROM3[905]<=26'd9774377; ROM4[905]<=26'd23487458;
ROM1[906]<=26'd2026704; ROM2[906]<=26'd11324226; ROM3[906]<=26'd9772467; ROM4[906]<=26'd23485537;
ROM1[907]<=26'd2039873; ROM2[907]<=26'd11328141; ROM3[907]<=26'd9770030; ROM4[907]<=26'd23487414;
ROM1[908]<=26'd2050496; ROM2[908]<=26'd11326291; ROM3[908]<=26'd9766027; ROM4[908]<=26'd23486197;
ROM1[909]<=26'd2047008; ROM2[909]<=26'd11324212; ROM3[909]<=26'd9765625; ROM4[909]<=26'd23485534;
ROM1[910]<=26'd2044988; ROM2[910]<=26'd11328209; ROM3[910]<=26'd9773233; ROM4[910]<=26'd23492195;
ROM1[911]<=26'd2042409; ROM2[911]<=26'd11331142; ROM3[911]<=26'd9782584; ROM4[911]<=26'd23496258;
ROM1[912]<=26'd2033111; ROM2[912]<=26'd11328785; ROM3[912]<=26'd9783769; ROM4[912]<=26'd23493421;
ROM1[913]<=26'd2021864; ROM2[913]<=26'd11324254; ROM3[913]<=26'd9783057; ROM4[913]<=26'd23489482;
ROM1[914]<=26'd2019824; ROM2[914]<=26'd11322521; ROM3[914]<=26'd9785367; ROM4[914]<=26'd23490795;
ROM1[915]<=26'd2025743; ROM2[915]<=26'd11322852; ROM3[915]<=26'd9786638; ROM4[915]<=26'd23494399;
ROM1[916]<=26'd2038083; ROM2[916]<=26'd11325327; ROM3[916]<=26'd9783230; ROM4[916]<=26'd23496071;
ROM1[917]<=26'd2045101; ROM2[917]<=26'd11328323; ROM3[917]<=26'd9781200; ROM4[917]<=26'd23497305;
ROM1[918]<=26'd2046146; ROM2[918]<=26'd11335279; ROM3[918]<=26'd9789583; ROM4[918]<=26'd23503621;
ROM1[919]<=26'd2026570; ROM2[919]<=26'd11322656; ROM3[919]<=26'd9781650; ROM4[919]<=26'd23493837;
ROM1[920]<=26'd2002761; ROM2[920]<=26'd11304623; ROM3[920]<=26'd9767671; ROM4[920]<=26'd23477503;
ROM1[921]<=26'd1994452; ROM2[921]<=26'd11304092; ROM3[921]<=26'd9771451; ROM4[921]<=26'd23477333;
ROM1[922]<=26'd1986695; ROM2[922]<=26'd11303299; ROM3[922]<=26'd9769904; ROM4[922]<=26'd23474827;
ROM1[923]<=26'd1996098; ROM2[923]<=26'd11310392; ROM3[923]<=26'd9770958; ROM4[923]<=26'd23476669;
ROM1[924]<=26'd2017970; ROM2[924]<=26'd11321967; ROM3[924]<=26'd9779117; ROM4[924]<=26'd23488015;
ROM1[925]<=26'd2021001; ROM2[925]<=26'd11317029; ROM3[925]<=26'd9771477; ROM4[925]<=26'd23485397;
ROM1[926]<=26'd2006564; ROM2[926]<=26'd11305811; ROM3[926]<=26'd9761939; ROM4[926]<=26'd23475596;
ROM1[927]<=26'd1999048; ROM2[927]<=26'd11308039; ROM3[927]<=26'd9767370; ROM4[927]<=26'd23478101;
ROM1[928]<=26'd1994682; ROM2[928]<=26'd11309545; ROM3[928]<=26'd9771783; ROM4[928]<=26'd23479689;
ROM1[929]<=26'd1978522; ROM2[929]<=26'd11299398; ROM3[929]<=26'd9764470; ROM4[929]<=26'd23470916;
ROM1[930]<=26'd1971853; ROM2[930]<=26'd11299512; ROM3[930]<=26'd9764372; ROM4[930]<=26'd23470032;
ROM1[931]<=26'd1970849; ROM2[931]<=26'd11298388; ROM3[931]<=26'd9763712; ROM4[931]<=26'd23470282;
ROM1[932]<=26'd1976709; ROM2[932]<=26'd11297047; ROM3[932]<=26'd9755738; ROM4[932]<=26'd23466466;
ROM1[933]<=26'd1993520; ROM2[933]<=26'd11304346; ROM3[933]<=26'd9750844; ROM4[933]<=26'd23468954;
ROM1[934]<=26'd1992591; ROM2[934]<=26'd11301820; ROM3[934]<=26'd9748129; ROM4[934]<=26'd23467371;
ROM1[935]<=26'd1982019; ROM2[935]<=26'd11297019; ROM3[935]<=26'd9747236; ROM4[935]<=26'd23464640;
ROM1[936]<=26'd1975754; ROM2[936]<=26'd11298601; ROM3[936]<=26'd9751728; ROM4[936]<=26'd23466784;
ROM1[937]<=26'd1971809; ROM2[937]<=26'd11299860; ROM3[937]<=26'd9759652; ROM4[937]<=26'd23471173;
ROM1[938]<=26'd1963523; ROM2[938]<=26'd11297800; ROM3[938]<=26'd9761426; ROM4[938]<=26'd23470400;
ROM1[939]<=26'd1961934; ROM2[939]<=26'd11299261; ROM3[939]<=26'd9760011; ROM4[939]<=26'd23467776;
ROM1[940]<=26'd1970344; ROM2[940]<=26'd11301511; ROM3[940]<=26'd9758061; ROM4[940]<=26'd23469376;
ROM1[941]<=26'd1984942; ROM2[941]<=26'd11305759; ROM3[941]<=26'd9754607; ROM4[941]<=26'd23471463;
ROM1[942]<=26'd1990443; ROM2[942]<=26'd11307219; ROM3[942]<=26'd9753769; ROM4[942]<=26'd23472848;
ROM1[943]<=26'd1988886; ROM2[943]<=26'd11309066; ROM3[943]<=26'd9760608; ROM4[943]<=26'd23477411;
ROM1[944]<=26'd1993563; ROM2[944]<=26'd11318875; ROM3[944]<=26'd9776250; ROM4[944]<=26'd23488322;
ROM1[945]<=26'd1985109; ROM2[945]<=26'd11315068; ROM3[945]<=26'd9777924; ROM4[945]<=26'd23485968;
ROM1[946]<=26'd1968525; ROM2[946]<=26'd11303069; ROM3[946]<=26'd9770624; ROM4[946]<=26'd23475613;
ROM1[947]<=26'd1959408; ROM2[947]<=26'd11295089; ROM3[947]<=26'd9764606; ROM4[947]<=26'd23469152;
ROM1[948]<=26'd1957017; ROM2[948]<=26'd11289954; ROM3[948]<=26'd9757571; ROM4[948]<=26'd23461786;
ROM1[949]<=26'd1973127; ROM2[949]<=26'd11294363; ROM3[949]<=26'd9757561; ROM4[949]<=26'd23465781;
ROM1[950]<=26'd1989328; ROM2[950]<=26'd11300879; ROM3[950]<=26'd9759264; ROM4[950]<=26'd23469925;
ROM1[951]<=26'd1986600; ROM2[951]<=26'd11301795; ROM3[951]<=26'd9760761; ROM4[951]<=26'd23469949;
ROM1[952]<=26'd1978099; ROM2[952]<=26'd11302801; ROM3[952]<=26'd9764431; ROM4[952]<=26'd23473325;
ROM1[953]<=26'd1982289; ROM2[953]<=26'd11314314; ROM3[953]<=26'd9775960; ROM4[953]<=26'd23483266;
ROM1[954]<=26'd1976247; ROM2[954]<=26'd11313843; ROM3[954]<=26'd9776470; ROM4[954]<=26'd23482454;
ROM1[955]<=26'd1960588; ROM2[955]<=26'd11301659; ROM3[955]<=26'd9767438; ROM4[955]<=26'd23470581;
ROM1[956]<=26'd1959614; ROM2[956]<=26'd11297823; ROM3[956]<=26'd9763674; ROM4[956]<=26'd23466571;
ROM1[957]<=26'd1959974; ROM2[957]<=26'd11290258; ROM3[957]<=26'd9752118; ROM4[957]<=26'd23456822;
ROM1[958]<=26'd1972771; ROM2[958]<=26'd11290646; ROM3[958]<=26'd9748658; ROM4[958]<=26'd23456741;
ROM1[959]<=26'd1980302; ROM2[959]<=26'd11296435; ROM3[959]<=26'd9754205; ROM4[959]<=26'd23462642;
ROM1[960]<=26'd1972429; ROM2[960]<=26'd11294539; ROM3[960]<=26'd9755053; ROM4[960]<=26'd23459711;
ROM1[961]<=26'd1969605; ROM2[961]<=26'd11296774; ROM3[961]<=26'd9762739; ROM4[961]<=26'd23462242;
ROM1[962]<=26'd1970992; ROM2[962]<=26'd11303626; ROM3[962]<=26'd9772469; ROM4[962]<=26'd23469152;
ROM1[963]<=26'd1968360; ROM2[963]<=26'd11305830; ROM3[963]<=26'd9776833; ROM4[963]<=26'd23472875;
ROM1[964]<=26'd1963957; ROM2[964]<=26'd11300985; ROM3[964]<=26'd9773473; ROM4[964]<=26'd23469613;
ROM1[965]<=26'd1966530; ROM2[965]<=26'd11296816; ROM3[965]<=26'd9767463; ROM4[965]<=26'd23466504;
ROM1[966]<=26'd1984669; ROM2[966]<=26'd11303110; ROM3[966]<=26'd9766719; ROM4[966]<=26'd23472187;
ROM1[967]<=26'd1990214; ROM2[967]<=26'd11304731; ROM3[967]<=26'd9764371; ROM4[967]<=26'd23473653;
ROM1[968]<=26'd1981520; ROM2[968]<=26'd11301103; ROM3[968]<=26'd9763069; ROM4[968]<=26'd23471428;
ROM1[969]<=26'd1975237; ROM2[969]<=26'd11299944; ROM3[969]<=26'd9767577; ROM4[969]<=26'd23472893;
ROM1[970]<=26'd1972138; ROM2[970]<=26'd11302055; ROM3[970]<=26'd9773853; ROM4[970]<=26'd23476054;
ROM1[971]<=26'd1970979; ROM2[971]<=26'd11304894; ROM3[971]<=26'd9779874; ROM4[971]<=26'd23479380;
ROM1[972]<=26'd1965858; ROM2[972]<=26'd11300872; ROM3[972]<=26'd9776616; ROM4[972]<=26'd23477213;
ROM1[973]<=26'd1968387; ROM2[973]<=26'd11301739; ROM3[973]<=26'd9773933; ROM4[973]<=26'd23477070;
ROM1[974]<=26'd1974483; ROM2[974]<=26'd11298858; ROM3[974]<=26'd9765555; ROM4[974]<=26'd23473293;
ROM1[975]<=26'd1976961; ROM2[975]<=26'd11294143; ROM3[975]<=26'd9755234; ROM4[975]<=26'd23467713;
ROM1[976]<=26'd1979442; ROM2[976]<=26'd11299953; ROM3[976]<=26'd9761335; ROM4[976]<=26'd23472880;
ROM1[977]<=26'd1971445; ROM2[977]<=26'd11297436; ROM3[977]<=26'd9762220; ROM4[977]<=26'd23471288;
ROM1[978]<=26'd1961070; ROM2[978]<=26'd11291990; ROM3[978]<=26'd9763081; ROM4[978]<=26'd23468314;
ROM1[979]<=26'd1957684; ROM2[979]<=26'd11294136; ROM3[979]<=26'd9770893; ROM4[979]<=26'd23472143;
ROM1[980]<=26'd1956613; ROM2[980]<=26'd11296832; ROM3[980]<=26'd9774971; ROM4[980]<=26'd23474366;
ROM1[981]<=26'd1957785; ROM2[981]<=26'd11298213; ROM3[981]<=26'd9772007; ROM4[981]<=26'd23472487;
ROM1[982]<=26'd1965009; ROM2[982]<=26'd11298580; ROM3[982]<=26'd9764550; ROM4[982]<=26'd23468678;
ROM1[983]<=26'd1978012; ROM2[983]<=26'd11301130; ROM3[983]<=26'd9760090; ROM4[983]<=26'd23470016;
ROM1[984]<=26'd1982812; ROM2[984]<=26'd11305404; ROM3[984]<=26'd9763476; ROM4[984]<=26'd23476209;
ROM1[985]<=26'd1974437; ROM2[985]<=26'd11302229; ROM3[985]<=26'd9764157; ROM4[985]<=26'd23476697;
ROM1[986]<=26'd1958245; ROM2[986]<=26'd11291660; ROM3[986]<=26'd9757055; ROM4[986]<=26'd23467080;
ROM1[987]<=26'd1955427; ROM2[987]<=26'd11293559; ROM3[987]<=26'd9760302; ROM4[987]<=26'd23469466;
ROM1[988]<=26'd1953819; ROM2[988]<=26'd11297167; ROM3[988]<=26'd9765253; ROM4[988]<=26'd23473677;
ROM1[989]<=26'd1952046; ROM2[989]<=26'd11295012; ROM3[989]<=26'd9762992; ROM4[989]<=26'd23470421;
ROM1[990]<=26'd1965601; ROM2[990]<=26'd11302723; ROM3[990]<=26'd9765274; ROM4[990]<=26'd23475066;
ROM1[991]<=26'd1978421; ROM2[991]<=26'd11305173; ROM3[991]<=26'd9759424; ROM4[991]<=26'd23474119;
ROM1[992]<=26'd1974824; ROM2[992]<=26'd11295226; ROM3[992]<=26'd9748120; ROM4[992]<=26'd23463949;
ROM1[993]<=26'd1973825; ROM2[993]<=26'd11298897; ROM3[993]<=26'd9753169; ROM4[993]<=26'd23467877;
ROM1[994]<=26'd1970673; ROM2[994]<=26'd11302627; ROM3[994]<=26'd9760952; ROM4[994]<=26'd23473036;
ROM1[995]<=26'd1958394; ROM2[995]<=26'd11294029; ROM3[995]<=26'd9758381; ROM4[995]<=26'd23466592;
ROM1[996]<=26'd1953335; ROM2[996]<=26'd11296363; ROM3[996]<=26'd9762537; ROM4[996]<=26'd23468297;
ROM1[997]<=26'd1950352; ROM2[997]<=26'd11296316; ROM3[997]<=26'd9763887; ROM4[997]<=26'd23467404;
ROM1[998]<=26'd1948887; ROM2[998]<=26'd11289468; ROM3[998]<=26'd9755493; ROM4[998]<=26'd23461485;
ROM1[999]<=26'd1960177; ROM2[999]<=26'd11291301; ROM3[999]<=26'd9752083; ROM4[999]<=26'd23461845;
ROM1[1000]<=26'd1966749; ROM2[1000]<=26'd11288817; ROM3[1000]<=26'd9747485; ROM4[1000]<=26'd23459951;
ROM1[1001]<=26'd1960831; ROM2[1001]<=26'd11283489; ROM3[1001]<=26'd9745973; ROM4[1001]<=26'd23458008;
ROM1[1002]<=26'd1954597; ROM2[1002]<=26'd11284556; ROM3[1002]<=26'd9753303; ROM4[1002]<=26'd23459464;
ROM1[1003]<=26'd1949537; ROM2[1003]<=26'd11286475; ROM3[1003]<=26'd9758535; ROM4[1003]<=26'd23460302;
ROM1[1004]<=26'd1943928; ROM2[1004]<=26'd11285044; ROM3[1004]<=26'd9758426; ROM4[1004]<=26'd23458267;
ROM1[1005]<=26'd1938401; ROM2[1005]<=26'd11283226; ROM3[1005]<=26'd9758392; ROM4[1005]<=26'd23456077;
ROM1[1006]<=26'd1941571; ROM2[1006]<=26'd11284069; ROM3[1006]<=26'd9757617; ROM4[1006]<=26'd23456693;
ROM1[1007]<=26'd1952092; ROM2[1007]<=26'd11284994; ROM3[1007]<=26'd9751069; ROM4[1007]<=26'd23455170;
ROM1[1008]<=26'd1964918; ROM2[1008]<=26'd11288596; ROM3[1008]<=26'd9746699; ROM4[1008]<=26'd23455245;
ROM1[1009]<=26'd1967563; ROM2[1009]<=26'd11290303; ROM3[1009]<=26'd9745376; ROM4[1009]<=26'd23456449;
ROM1[1010]<=26'd1962318; ROM2[1010]<=26'd11292124; ROM3[1010]<=26'd9746666; ROM4[1010]<=26'd23457641;
ROM1[1011]<=26'd1957341; ROM2[1011]<=26'd11293194; ROM3[1011]<=26'd9752196; ROM4[1011]<=26'd23460035;
ROM1[1012]<=26'd1952705; ROM2[1012]<=26'd11293217; ROM3[1012]<=26'd9756499; ROM4[1012]<=26'd23463014;
ROM1[1013]<=26'd1949663; ROM2[1013]<=26'd11296117; ROM3[1013]<=26'd9761458; ROM4[1013]<=26'd23465692;
ROM1[1014]<=26'd1955939; ROM2[1014]<=26'd11300995; ROM3[1014]<=26'd9766873; ROM4[1014]<=26'd23472062;
ROM1[1015]<=26'd1968646; ROM2[1015]<=26'd11305768; ROM3[1015]<=26'd9768085; ROM4[1015]<=26'd23476625;
ROM1[1016]<=26'd1980042; ROM2[1016]<=26'd11305354; ROM3[1016]<=26'd9763698; ROM4[1016]<=26'd23474944;
ROM1[1017]<=26'd1983366; ROM2[1017]<=26'd11304639; ROM3[1017]<=26'd9760993; ROM4[1017]<=26'd23474510;
ROM1[1018]<=26'd1981781; ROM2[1018]<=26'd11307336; ROM3[1018]<=26'd9766506; ROM4[1018]<=26'd23478015;
ROM1[1019]<=26'd1977832; ROM2[1019]<=26'd11310377; ROM3[1019]<=26'd9774018; ROM4[1019]<=26'd23482234;
ROM1[1020]<=26'd1966634; ROM2[1020]<=26'd11305637; ROM3[1020]<=26'd9771215; ROM4[1020]<=26'd23477432;
ROM1[1021]<=26'd1955976; ROM2[1021]<=26'd11300350; ROM3[1021]<=26'd9769308; ROM4[1021]<=26'd23473232;
ROM1[1022]<=26'd1956816; ROM2[1022]<=26'd11303350; ROM3[1022]<=26'd9771029; ROM4[1022]<=26'd23474686;
ROM1[1023]<=26'd1962278; ROM2[1023]<=26'd11304142; ROM3[1023]<=26'd9767639; ROM4[1023]<=26'd23473458;
ROM1[1024]<=26'd1975285; ROM2[1024]<=26'd11304230; ROM3[1024]<=26'd9763072; ROM4[1024]<=26'd23471398;
ROM1[1025]<=26'd1984997; ROM2[1025]<=26'd11305019; ROM3[1025]<=26'd9759493; ROM4[1025]<=26'd23471997;
ROM1[1026]<=26'd1972198; ROM2[1026]<=26'd11295298; ROM3[1026]<=26'd9752980; ROM4[1026]<=26'd23464297;
ROM1[1027]<=26'd1958762; ROM2[1027]<=26'd11289916; ROM3[1027]<=26'd9751128; ROM4[1027]<=26'd23458296;
ROM1[1028]<=26'd1957980; ROM2[1028]<=26'd11295634; ROM3[1028]<=26'd9756973; ROM4[1028]<=26'd23464822;
ROM1[1029]<=26'd1956407; ROM2[1029]<=26'd11298726; ROM3[1029]<=26'd9762368; ROM4[1029]<=26'd23469227;
ROM1[1030]<=26'd1954244; ROM2[1030]<=26'd11298670; ROM3[1030]<=26'd9763344; ROM4[1030]<=26'd23469848;
ROM1[1031]<=26'd1956086; ROM2[1031]<=26'd11296794; ROM3[1031]<=26'd9760069; ROM4[1031]<=26'd23468522;
ROM1[1032]<=26'd1963353; ROM2[1032]<=26'd11294446; ROM3[1032]<=26'd9753330; ROM4[1032]<=26'd23465704;
ROM1[1033]<=26'd1972779; ROM2[1033]<=26'd11292764; ROM3[1033]<=26'd9745089; ROM4[1033]<=26'd23463635;
ROM1[1034]<=26'd1975430; ROM2[1034]<=26'd11294434; ROM3[1034]<=26'd9745058; ROM4[1034]<=26'd23464750;
ROM1[1035]<=26'd1967731; ROM2[1035]<=26'd11292940; ROM3[1035]<=26'd9745265; ROM4[1035]<=26'd23464500;
ROM1[1036]<=26'd1959010; ROM2[1036]<=26'd11289832; ROM3[1036]<=26'd9746410; ROM4[1036]<=26'd23462081;
ROM1[1037]<=26'd1956565; ROM2[1037]<=26'd11294256; ROM3[1037]<=26'd9751346; ROM4[1037]<=26'd23464568;
ROM1[1038]<=26'd1954089; ROM2[1038]<=26'd11298832; ROM3[1038]<=26'd9757236; ROM4[1038]<=26'd23470629;
ROM1[1039]<=26'd1954308; ROM2[1039]<=26'd11298723; ROM3[1039]<=26'd9758620; ROM4[1039]<=26'd23470694;
ROM1[1040]<=26'd1962249; ROM2[1040]<=26'd11300811; ROM3[1040]<=26'd9756906; ROM4[1040]<=26'd23471124;
ROM1[1041]<=26'd1971210; ROM2[1041]<=26'd11298596; ROM3[1041]<=26'd9749623; ROM4[1041]<=26'd23467389;
ROM1[1042]<=26'd1969479; ROM2[1042]<=26'd11291426; ROM3[1042]<=26'd9742216; ROM4[1042]<=26'd23459563;
ROM1[1043]<=26'd1967550; ROM2[1043]<=26'd11293745; ROM3[1043]<=26'd9748051; ROM4[1043]<=26'd23464478;
ROM1[1044]<=26'd1960843; ROM2[1044]<=26'd11293433; ROM3[1044]<=26'd9751908; ROM4[1044]<=26'd23465477;
ROM1[1045]<=26'd1954991; ROM2[1045]<=26'd11291909; ROM3[1045]<=26'd9753489; ROM4[1045]<=26'd23465610;
ROM1[1046]<=26'd1949841; ROM2[1046]<=26'd11291626; ROM3[1046]<=26'd9756687; ROM4[1046]<=26'd23466751;
ROM1[1047]<=26'd1945235; ROM2[1047]<=26'd11288565; ROM3[1047]<=26'd9756026; ROM4[1047]<=26'd23463340;
ROM1[1048]<=26'd1950077; ROM2[1048]<=26'd11289470; ROM3[1048]<=26'd9754405; ROM4[1048]<=26'd23463648;
ROM1[1049]<=26'd1963184; ROM2[1049]<=26'd11292074; ROM3[1049]<=26'd9750070; ROM4[1049]<=26'd23463600;
ROM1[1050]<=26'd1971131; ROM2[1050]<=26'd11292492; ROM3[1050]<=26'd9746114; ROM4[1050]<=26'd23462632;
ROM1[1051]<=26'd1965779; ROM2[1051]<=26'd11292252; ROM3[1051]<=26'd9746448; ROM4[1051]<=26'd23461789;
ROM1[1052]<=26'd1962350; ROM2[1052]<=26'd11297650; ROM3[1052]<=26'd9756150; ROM4[1052]<=26'd23466978;
ROM1[1053]<=26'd1959946; ROM2[1053]<=26'd11300159; ROM3[1053]<=26'd9764153; ROM4[1053]<=26'd23470174;
ROM1[1054]<=26'd1951427; ROM2[1054]<=26'd11296304; ROM3[1054]<=26'd9762601; ROM4[1054]<=26'd23466749;
ROM1[1055]<=26'd1953021; ROM2[1055]<=26'd11300349; ROM3[1055]<=26'd9767136; ROM4[1055]<=26'd23470584;
ROM1[1056]<=26'd1961251; ROM2[1056]<=26'd11305764; ROM3[1056]<=26'd9770552; ROM4[1056]<=26'd23475977;
ROM1[1057]<=26'd1964088; ROM2[1057]<=26'd11300418; ROM3[1057]<=26'd9761110; ROM4[1057]<=26'd23469724;
ROM1[1058]<=26'd1972335; ROM2[1058]<=26'd11296808; ROM3[1058]<=26'd9752297; ROM4[1058]<=26'd23464992;
ROM1[1059]<=26'd1974340; ROM2[1059]<=26'd11298229; ROM3[1059]<=26'd9753906; ROM4[1059]<=26'd23467731;
ROM1[1060]<=26'd1964402; ROM2[1060]<=26'd11292409; ROM3[1060]<=26'd9752007; ROM4[1060]<=26'd23464057;
ROM1[1061]<=26'd1958414; ROM2[1061]<=26'd11292880; ROM3[1061]<=26'd9757493; ROM4[1061]<=26'd23465890;
ROM1[1062]<=26'd1953512; ROM2[1062]<=26'd11295631; ROM3[1062]<=26'd9761053; ROM4[1062]<=26'd23468424;
ROM1[1063]<=26'd1945340; ROM2[1063]<=26'd11293439; ROM3[1063]<=26'd9758973; ROM4[1063]<=26'd23464509;
ROM1[1064]<=26'd1945564; ROM2[1064]<=26'd11293516; ROM3[1064]<=26'd9758081; ROM4[1064]<=26'd23462986;
ROM1[1065]<=26'd1950995; ROM2[1065]<=26'd11292078; ROM3[1065]<=26'd9750608; ROM4[1065]<=26'd23460263;
ROM1[1066]<=26'd1963408; ROM2[1066]<=26'd11293808; ROM3[1066]<=26'd9746850; ROM4[1066]<=26'd23459294;
ROM1[1067]<=26'd1964460; ROM2[1067]<=26'd11292860; ROM3[1067]<=26'd9743201; ROM4[1067]<=26'd23456222;
ROM1[1068]<=26'd1956843; ROM2[1068]<=26'd11290164; ROM3[1068]<=26'd9740535; ROM4[1068]<=26'd23454133;
ROM1[1069]<=26'd1952807; ROM2[1069]<=26'd11292605; ROM3[1069]<=26'd9746711; ROM4[1069]<=26'd23457944;
ROM1[1070]<=26'd1950379; ROM2[1070]<=26'd11296966; ROM3[1070]<=26'd9754815; ROM4[1070]<=26'd23462395;
ROM1[1071]<=26'd1945465; ROM2[1071]<=26'd11295987; ROM3[1071]<=26'd9759145; ROM4[1071]<=26'd23464574;
ROM1[1072]<=26'd1940740; ROM2[1072]<=26'd11294710; ROM3[1072]<=26'd9758462; ROM4[1072]<=26'd23462091;
ROM1[1073]<=26'd1949806; ROM2[1073]<=26'd11300086; ROM3[1073]<=26'd9760848; ROM4[1073]<=26'd23465497;
ROM1[1074]<=26'd1971873; ROM2[1074]<=26'd11309233; ROM3[1074]<=26'd9763831; ROM4[1074]<=26'd23474459;
ROM1[1075]<=26'd1975078; ROM2[1075]<=26'd11304060; ROM3[1075]<=26'd9751361; ROM4[1075]<=26'd23468184;
ROM1[1076]<=26'd1960098; ROM2[1076]<=26'd11291862; ROM3[1076]<=26'd9741143; ROM4[1076]<=26'd23456720;
ROM1[1077]<=26'd1950048; ROM2[1077]<=26'd11287450; ROM3[1077]<=26'd9741026; ROM4[1077]<=26'd23453160;
ROM1[1078]<=26'd1939541; ROM2[1078]<=26'd11281329; ROM3[1078]<=26'd9740205; ROM4[1078]<=26'd23449576;
ROM1[1079]<=26'd1937037; ROM2[1079]<=26'd11283473; ROM3[1079]<=26'd9746842; ROM4[1079]<=26'd23453720;
ROM1[1080]<=26'd1943032; ROM2[1080]<=26'd11293195; ROM3[1080]<=26'd9757207; ROM4[1080]<=26'd23465863;
ROM1[1081]<=26'd1949585; ROM2[1081]<=26'd11297728; ROM3[1081]<=26'd9759083; ROM4[1081]<=26'd23470463;
ROM1[1082]<=26'd1956232; ROM2[1082]<=26'd11296599; ROM3[1082]<=26'd9750571; ROM4[1082]<=26'd23464104;
ROM1[1083]<=26'd1966831; ROM2[1083]<=26'd11297104; ROM3[1083]<=26'd9744257; ROM4[1083]<=26'd23462697;
ROM1[1084]<=26'd1967233; ROM2[1084]<=26'd11296130; ROM3[1084]<=26'd9743920; ROM4[1084]<=26'd23462519;
ROM1[1085]<=26'd1959880; ROM2[1085]<=26'd11293736; ROM3[1085]<=26'd9745919; ROM4[1085]<=26'd23460968;
ROM1[1086]<=26'd1959116; ROM2[1086]<=26'd11297856; ROM3[1086]<=26'd9754248; ROM4[1086]<=26'd23467926;
ROM1[1087]<=26'd1949944; ROM2[1087]<=26'd11292598; ROM3[1087]<=26'd9752862; ROM4[1087]<=26'd23464027;
ROM1[1088]<=26'd1937378; ROM2[1088]<=26'd11284134; ROM3[1088]<=26'd9748795; ROM4[1088]<=26'd23455064;
ROM1[1089]<=26'd1936607; ROM2[1089]<=26'd11283638; ROM3[1089]<=26'd9749592; ROM4[1089]<=26'd23453167;
ROM1[1090]<=26'd1947947; ROM2[1090]<=26'd11288084; ROM3[1090]<=26'd9750772; ROM4[1090]<=26'd23456904;
ROM1[1091]<=26'd1965554; ROM2[1091]<=26'd11293747; ROM3[1091]<=26'd9749443; ROM4[1091]<=26'd23461968;
ROM1[1092]<=26'd1967740; ROM2[1092]<=26'd11290544; ROM3[1092]<=26'd9742438; ROM4[1092]<=26'd23457554;
ROM1[1093]<=26'd1959080; ROM2[1093]<=26'd11287962; ROM3[1093]<=26'd9744420; ROM4[1093]<=26'd23456414;
ROM1[1094]<=26'd1945169; ROM2[1094]<=26'd11283620; ROM3[1094]<=26'd9745151; ROM4[1094]<=26'd23452751;
ROM1[1095]<=26'd1937852; ROM2[1095]<=26'd11280966; ROM3[1095]<=26'd9748038; ROM4[1095]<=26'd23451400;
ROM1[1096]<=26'd1937024; ROM2[1096]<=26'd11284911; ROM3[1096]<=26'd9757358; ROM4[1096]<=26'd23457911;
ROM1[1097]<=26'd1937860; ROM2[1097]<=26'd11286668; ROM3[1097]<=26'd9758736; ROM4[1097]<=26'd23459144;
ROM1[1098]<=26'd1941454; ROM2[1098]<=26'd11284852; ROM3[1098]<=26'd9753714; ROM4[1098]<=26'd23457955;
ROM1[1099]<=26'd1955883; ROM2[1099]<=26'd11287925; ROM3[1099]<=26'd9750520; ROM4[1099]<=26'd23459941;
ROM1[1100]<=26'd1966937; ROM2[1100]<=26'd11290599; ROM3[1100]<=26'd9747404; ROM4[1100]<=26'd23460834;
ROM1[1101]<=26'd1961090; ROM2[1101]<=26'd11288492; ROM3[1101]<=26'd9744764; ROM4[1101]<=26'd23459851;
ROM1[1102]<=26'd1953014; ROM2[1102]<=26'd11285709; ROM3[1102]<=26'd9748985; ROM4[1102]<=26'd23459865;
ROM1[1103]<=26'd1948898; ROM2[1103]<=26'd11286845; ROM3[1103]<=26'd9755807; ROM4[1103]<=26'd23462384;
ROM1[1104]<=26'd1949294; ROM2[1104]<=26'd11292981; ROM3[1104]<=26'd9765804; ROM4[1104]<=26'd23470130;
ROM1[1105]<=26'd1948689; ROM2[1105]<=26'd11294099; ROM3[1105]<=26'd9771409; ROM4[1105]<=26'd23473009;
ROM1[1106]<=26'd1949175; ROM2[1106]<=26'd11292198; ROM3[1106]<=26'd9765709; ROM4[1106]<=26'd23469674;
ROM1[1107]<=26'd1959323; ROM2[1107]<=26'd11292634; ROM3[1107]<=26'd9760122; ROM4[1107]<=26'd23468176;
ROM1[1108]<=26'd1974841; ROM2[1108]<=26'd11296776; ROM3[1108]<=26'd9760240; ROM4[1108]<=26'd23470201;
ROM1[1109]<=26'd1972389; ROM2[1109]<=26'd11293013; ROM3[1109]<=26'd9755850; ROM4[1109]<=26'd23466123;
ROM1[1110]<=26'd1962278; ROM2[1110]<=26'd11288204; ROM3[1110]<=26'd9755877; ROM4[1110]<=26'd23462910;
ROM1[1111]<=26'd1955575; ROM2[1111]<=26'd11288442; ROM3[1111]<=26'd9761541; ROM4[1111]<=26'd23464629;
ROM1[1112]<=26'd1949111; ROM2[1112]<=26'd11289262; ROM3[1112]<=26'd9762623; ROM4[1112]<=26'd23464904;
ROM1[1113]<=26'd1942006; ROM2[1113]<=26'd11287081; ROM3[1113]<=26'd9764639; ROM4[1113]<=26'd23464885;
ROM1[1114]<=26'd1936343; ROM2[1114]<=26'd11282403; ROM3[1114]<=26'd9758966; ROM4[1114]<=26'd23459555;
ROM1[1115]<=26'd1939903; ROM2[1115]<=26'd11281523; ROM3[1115]<=26'd9752977; ROM4[1115]<=26'd23456453;
ROM1[1116]<=26'd1952241; ROM2[1116]<=26'd11281814; ROM3[1116]<=26'd9749071; ROM4[1116]<=26'd23456298;
ROM1[1117]<=26'd1964204; ROM2[1117]<=26'd11289976; ROM3[1117]<=26'd9751790; ROM4[1117]<=26'd23462130;
ROM1[1118]<=26'd1969473; ROM2[1118]<=26'd11298526; ROM3[1118]<=26'd9762936; ROM4[1118]<=26'd23472438;
ROM1[1119]<=26'd1957183; ROM2[1119]<=26'd11292430; ROM3[1119]<=26'd9760855; ROM4[1119]<=26'd23467547;
ROM1[1120]<=26'd1943891; ROM2[1120]<=26'd11284904; ROM3[1120]<=26'd9755816; ROM4[1120]<=26'd23462588;
ROM1[1121]<=26'd1938777; ROM2[1121]<=26'd11283455; ROM3[1121]<=26'd9759157; ROM4[1121]<=26'd23462443;
ROM1[1122]<=26'd1939046; ROM2[1122]<=26'd11285513; ROM3[1122]<=26'd9760225; ROM4[1122]<=26'd23462744;
ROM1[1123]<=26'd1949375; ROM2[1123]<=26'd11289781; ROM3[1123]<=26'd9760690; ROM4[1123]<=26'd23465632;
ROM1[1124]<=26'd1962845; ROM2[1124]<=26'd11293472; ROM3[1124]<=26'd9759588; ROM4[1124]<=26'd23467735;
ROM1[1125]<=26'd1971769; ROM2[1125]<=26'd11298030; ROM3[1125]<=26'd9755934; ROM4[1125]<=26'd23470523;
ROM1[1126]<=26'd1966814; ROM2[1126]<=26'd11294904; ROM3[1126]<=26'd9752062; ROM4[1126]<=26'd23466165;
ROM1[1127]<=26'd1954341; ROM2[1127]<=26'd11288940; ROM3[1127]<=26'd9748552; ROM4[1127]<=26'd23461075;
ROM1[1128]<=26'd1947379; ROM2[1128]<=26'd11286594; ROM3[1128]<=26'd9747819; ROM4[1128]<=26'd23458925;
ROM1[1129]<=26'd1939347; ROM2[1129]<=26'd11282421; ROM3[1129]<=26'd9747916; ROM4[1129]<=26'd23455869;
ROM1[1130]<=26'd1936127; ROM2[1130]<=26'd11283759; ROM3[1130]<=26'd9750730; ROM4[1130]<=26'd23457362;
ROM1[1131]<=26'd1943064; ROM2[1131]<=26'd11289518; ROM3[1131]<=26'd9753709; ROM4[1131]<=26'd23460837;
ROM1[1132]<=26'd1955597; ROM2[1132]<=26'd11294405; ROM3[1132]<=26'd9753009; ROM4[1132]<=26'd23462974;
ROM1[1133]<=26'd1966266; ROM2[1133]<=26'd11294406; ROM3[1133]<=26'd9747505; ROM4[1133]<=26'd23462616;
ROM1[1134]<=26'd1965886; ROM2[1134]<=26'd11294321; ROM3[1134]<=26'd9746946; ROM4[1134]<=26'd23462531;
ROM1[1135]<=26'd1967106; ROM2[1135]<=26'd11301174; ROM3[1135]<=26'd9757184; ROM4[1135]<=26'd23470789;
ROM1[1136]<=26'd1962159; ROM2[1136]<=26'd11301990; ROM3[1136]<=26'd9763926; ROM4[1136]<=26'd23474013;
ROM1[1137]<=26'd1950709; ROM2[1137]<=26'd11295855; ROM3[1137]<=26'd9760033; ROM4[1137]<=26'd23467663;
ROM1[1138]<=26'd1942822; ROM2[1138]<=26'd11292102; ROM3[1138]<=26'd9757335; ROM4[1138]<=26'd23465304;
ROM1[1139]<=26'd1938167; ROM2[1139]<=26'd11288123; ROM3[1139]<=26'd9754420; ROM4[1139]<=26'd23462284;
ROM1[1140]<=26'd1942879; ROM2[1140]<=26'd11282434; ROM3[1140]<=26'd9747740; ROM4[1140]<=26'd23457790;
ROM1[1141]<=26'd1957248; ROM2[1141]<=26'd11284011; ROM3[1141]<=26'd9743854; ROM4[1141]<=26'd23459607;
ROM1[1142]<=26'd1962335; ROM2[1142]<=26'd11285619; ROM3[1142]<=26'd9745888; ROM4[1142]<=26'd23461160;
ROM1[1143]<=26'd1957428; ROM2[1143]<=26'd11282841; ROM3[1143]<=26'd9748423; ROM4[1143]<=26'd23460402;
ROM1[1144]<=26'd1952104; ROM2[1144]<=26'd11286703; ROM3[1144]<=26'd9755079; ROM4[1144]<=26'd23464762;
ROM1[1145]<=26'd1949071; ROM2[1145]<=26'd11290524; ROM3[1145]<=26'd9763509; ROM4[1145]<=26'd23469992;
ROM1[1146]<=26'd1940741; ROM2[1146]<=26'd11288465; ROM3[1146]<=26'd9766451; ROM4[1146]<=26'd23470762;
ROM1[1147]<=26'd1938145; ROM2[1147]<=26'd11287618; ROM3[1147]<=26'd9767943; ROM4[1147]<=26'd23470563;
ROM1[1148]<=26'd1942823; ROM2[1148]<=26'd11287962; ROM3[1148]<=26'd9764989; ROM4[1148]<=26'd23468832;
ROM1[1149]<=26'd1955071; ROM2[1149]<=26'd11289214; ROM3[1149]<=26'd9759168; ROM4[1149]<=26'd23468358;
ROM1[1150]<=26'd1967673; ROM2[1150]<=26'd11293447; ROM3[1150]<=26'd9758789; ROM4[1150]<=26'd23472150;
ROM1[1151]<=26'd1965511; ROM2[1151]<=26'd11293870; ROM3[1151]<=26'd9759461; ROM4[1151]<=26'd23473147;
ROM1[1152]<=26'd1957270; ROM2[1152]<=26'd11291456; ROM3[1152]<=26'd9759555; ROM4[1152]<=26'd23470538;
ROM1[1153]<=26'd1950909; ROM2[1153]<=26'd11290830; ROM3[1153]<=26'd9760958; ROM4[1153]<=26'd23468485;
ROM1[1154]<=26'd1945023; ROM2[1154]<=26'd11290061; ROM3[1154]<=26'd9761539; ROM4[1154]<=26'd23465813;
ROM1[1155]<=26'd1940531; ROM2[1155]<=26'd11291532; ROM3[1155]<=26'd9761940; ROM4[1155]<=26'd23465522;
ROM1[1156]<=26'd1946034; ROM2[1156]<=26'd11294992; ROM3[1156]<=26'd9762917; ROM4[1156]<=26'd23468870;
ROM1[1157]<=26'd1958088; ROM2[1157]<=26'd11297522; ROM3[1157]<=26'd9761807; ROM4[1157]<=26'd23470843;
ROM1[1158]<=26'd1968812; ROM2[1158]<=26'd11298720; ROM3[1158]<=26'd9758522; ROM4[1158]<=26'd23470538;
ROM1[1159]<=26'd1971550; ROM2[1159]<=26'd11300091; ROM3[1159]<=26'd9759531; ROM4[1159]<=26'd23471918;
ROM1[1160]<=26'd1970619; ROM2[1160]<=26'd11302237; ROM3[1160]<=26'd9766561; ROM4[1160]<=26'd23478002;
ROM1[1161]<=26'd1960330; ROM2[1161]<=26'd11297273; ROM3[1161]<=26'd9767443; ROM4[1161]<=26'd23476170;
ROM1[1162]<=26'd1949182; ROM2[1162]<=26'd11290205; ROM3[1162]<=26'd9764225; ROM4[1162]<=26'd23471101;
ROM1[1163]<=26'd1944428; ROM2[1163]<=26'd11291263; ROM3[1163]<=26'd9768783; ROM4[1163]<=26'd23472870;
ROM1[1164]<=26'd1944353; ROM2[1164]<=26'd11291462; ROM3[1164]<=26'd9768373; ROM4[1164]<=26'd23471698;
ROM1[1165]<=26'd1953736; ROM2[1165]<=26'd11294899; ROM3[1165]<=26'd9766780; ROM4[1165]<=26'd23473734;
ROM1[1166]<=26'd1971848; ROM2[1166]<=26'd11301993; ROM3[1166]<=26'd9768322; ROM4[1166]<=26'd23478789;
ROM1[1167]<=26'd1976137; ROM2[1167]<=26'd11301445; ROM3[1167]<=26'd9765143; ROM4[1167]<=26'd23478806;
ROM1[1168]<=26'd1964913; ROM2[1168]<=26'd11294922; ROM3[1168]<=26'd9760885; ROM4[1168]<=26'd23473073;
ROM1[1169]<=26'd1955283; ROM2[1169]<=26'd11291813; ROM3[1169]<=26'd9761918; ROM4[1169]<=26'd23469509;
ROM1[1170]<=26'd1949408; ROM2[1170]<=26'd11291392; ROM3[1170]<=26'd9762515; ROM4[1170]<=26'd23469013;
ROM1[1171]<=26'd1943581; ROM2[1171]<=26'd11289920; ROM3[1171]<=26'd9764993; ROM4[1171]<=26'd23468459;
ROM1[1172]<=26'd1944167; ROM2[1172]<=26'd11294618; ROM3[1172]<=26'd9768409; ROM4[1172]<=26'd23471522;
ROM1[1173]<=26'd1949476; ROM2[1173]<=26'd11296104; ROM3[1173]<=26'd9766145; ROM4[1173]<=26'd23470723;
ROM1[1174]<=26'd1962052; ROM2[1174]<=26'd11295198; ROM3[1174]<=26'd9760530; ROM4[1174]<=26'd23470619;
ROM1[1175]<=26'd1971351; ROM2[1175]<=26'd11297598; ROM3[1175]<=26'd9757851; ROM4[1175]<=26'd23472168;
ROM1[1176]<=26'd1966249; ROM2[1176]<=26'd11295283; ROM3[1176]<=26'd9758586; ROM4[1176]<=26'd23470762;
ROM1[1177]<=26'd1959733; ROM2[1177]<=26'd11294487; ROM3[1177]<=26'd9760608; ROM4[1177]<=26'd23472336;
ROM1[1178]<=26'd1957110; ROM2[1178]<=26'd11298676; ROM3[1178]<=26'd9766203; ROM4[1178]<=26'd23476595;
ROM1[1179]<=26'd1959190; ROM2[1179]<=26'd11306104; ROM3[1179]<=26'd9775288; ROM4[1179]<=26'd23483267;
ROM1[1180]<=26'd1953218; ROM2[1180]<=26'd11304361; ROM3[1180]<=26'd9773040; ROM4[1180]<=26'd23480048;
ROM1[1181]<=26'd1943608; ROM2[1181]<=26'd11291365; ROM3[1181]<=26'd9759924; ROM4[1181]<=26'd23467109;
ROM1[1182]<=26'd1949582; ROM2[1182]<=26'd11287523; ROM3[1182]<=26'd9750943; ROM4[1182]<=26'd23461042;
ROM1[1183]<=26'd1956118; ROM2[1183]<=26'd11284605; ROM3[1183]<=26'd9742108; ROM4[1183]<=26'd23456498;
ROM1[1184]<=26'd1956035; ROM2[1184]<=26'd11285207; ROM3[1184]<=26'd9743267; ROM4[1184]<=26'd23457839;
ROM1[1185]<=26'd1957412; ROM2[1185]<=26'd11293372; ROM3[1185]<=26'd9752971; ROM4[1185]<=26'd23466747;
ROM1[1186]<=26'd1948586; ROM2[1186]<=26'd11291048; ROM3[1186]<=26'd9756245; ROM4[1186]<=26'd23464586;
ROM1[1187]<=26'd1937015; ROM2[1187]<=26'd11282489; ROM3[1187]<=26'd9750100; ROM4[1187]<=26'd23456869;
ROM1[1188]<=26'd1932735; ROM2[1188]<=26'd11281837; ROM3[1188]<=26'd9750075; ROM4[1188]<=26'd23456615;
ROM1[1189]<=26'd1939141; ROM2[1189]<=26'd11286982; ROM3[1189]<=26'd9754787; ROM4[1189]<=26'd23459978;
ROM1[1190]<=26'd1948466; ROM2[1190]<=26'd11288388; ROM3[1190]<=26'd9751017; ROM4[1190]<=26'd23460051;
ROM1[1191]<=26'd1960992; ROM2[1191]<=26'd11289530; ROM3[1191]<=26'd9747778; ROM4[1191]<=26'd23460416;
ROM1[1192]<=26'd1971264; ROM2[1192]<=26'd11295440; ROM3[1192]<=26'd9754367; ROM4[1192]<=26'd23466258;
ROM1[1193]<=26'd1976322; ROM2[1193]<=26'd11307327; ROM3[1193]<=26'd9767545; ROM4[1193]<=26'd23477520;
ROM1[1194]<=26'd1963050; ROM2[1194]<=26'd11301333; ROM3[1194]<=26'd9764798; ROM4[1194]<=26'd23473160;
ROM1[1195]<=26'd1948106; ROM2[1195]<=26'd11290142; ROM3[1195]<=26'd9757109; ROM4[1195]<=26'd23462784;
ROM1[1196]<=26'd1939447; ROM2[1196]<=26'd11287205; ROM3[1196]<=26'd9755897; ROM4[1196]<=26'd23459805;
ROM1[1197]<=26'd1935886; ROM2[1197]<=26'd11282938; ROM3[1197]<=26'd9753863; ROM4[1197]<=26'd23456520;
ROM1[1198]<=26'd1949917; ROM2[1198]<=26'd11288270; ROM3[1198]<=26'd9759604; ROM4[1198]<=26'd23463607;
ROM1[1199]<=26'd1973748; ROM2[1199]<=26'd11300359; ROM3[1199]<=26'd9766947; ROM4[1199]<=26'd23475301;
ROM1[1200]<=26'd1987425; ROM2[1200]<=26'd11304890; ROM3[1200]<=26'd9768673; ROM4[1200]<=26'd23480642;
ROM1[1201]<=26'd1976123; ROM2[1201]<=26'd11297225; ROM3[1201]<=26'd9763628; ROM4[1201]<=26'd23474686;
ROM1[1202]<=26'd1963321; ROM2[1202]<=26'd11292690; ROM3[1202]<=26'd9760592; ROM4[1202]<=26'd23469610;
ROM1[1203]<=26'd1955904; ROM2[1203]<=26'd11290463; ROM3[1203]<=26'd9762564; ROM4[1203]<=26'd23470597;
ROM1[1204]<=26'd1947942; ROM2[1204]<=26'd11288895; ROM3[1204]<=26'd9763412; ROM4[1204]<=26'd23469417;
ROM1[1205]<=26'd1949564; ROM2[1205]<=26'd11293300; ROM3[1205]<=26'd9768110; ROM4[1205]<=26'd23471565;
ROM1[1206]<=26'd1955951; ROM2[1206]<=26'd11294018; ROM3[1206]<=26'd9767854; ROM4[1206]<=26'd23472016;
ROM1[1207]<=26'd1960525; ROM2[1207]<=26'd11289833; ROM3[1207]<=26'd9755951; ROM4[1207]<=26'd23464980;
ROM1[1208]<=26'd1968566; ROM2[1208]<=26'd11286893; ROM3[1208]<=26'd9749347; ROM4[1208]<=26'd23462230;
ROM1[1209]<=26'd1966712; ROM2[1209]<=26'd11284644; ROM3[1209]<=26'd9748910; ROM4[1209]<=26'd23461532;
ROM1[1210]<=26'd1961603; ROM2[1210]<=26'd11288924; ROM3[1210]<=26'd9756139; ROM4[1210]<=26'd23465502;
ROM1[1211]<=26'd1956834; ROM2[1211]<=26'd11291378; ROM3[1211]<=26'd9762850; ROM4[1211]<=26'd23468306;
ROM1[1212]<=26'd1945899; ROM2[1212]<=26'd11285198; ROM3[1212]<=26'd9757487; ROM4[1212]<=26'd23462368;
ROM1[1213]<=26'd1935809; ROM2[1213]<=26'd11280521; ROM3[1213]<=26'd9754742; ROM4[1213]<=26'd23458317;
ROM1[1214]<=26'd1940010; ROM2[1214]<=26'd11283523; ROM3[1214]<=26'd9757324; ROM4[1214]<=26'd23461070;
ROM1[1215]<=26'd1956228; ROM2[1215]<=26'd11292462; ROM3[1215]<=26'd9761277; ROM4[1215]<=26'd23467404;
ROM1[1216]<=26'd1969487; ROM2[1216]<=26'd11293159; ROM3[1216]<=26'd9758251; ROM4[1216]<=26'd23468248;
ROM1[1217]<=26'd1967451; ROM2[1217]<=26'd11286994; ROM3[1217]<=26'd9751345; ROM4[1217]<=26'd23463921;
ROM1[1218]<=26'd1964090; ROM2[1218]<=26'd11289992; ROM3[1218]<=26'd9756832; ROM4[1218]<=26'd23467694;
ROM1[1219]<=26'd1960635; ROM2[1219]<=26'd11293987; ROM3[1219]<=26'd9764072; ROM4[1219]<=26'd23472974;
ROM1[1220]<=26'd1952192; ROM2[1220]<=26'd11288982; ROM3[1220]<=26'd9760558; ROM4[1220]<=26'd23468539;
ROM1[1221]<=26'd1942494; ROM2[1221]<=26'd11283060; ROM3[1221]<=26'd9758393; ROM4[1221]<=26'd23465035;
ROM1[1222]<=26'd1938408; ROM2[1222]<=26'd11280913; ROM3[1222]<=26'd9756454; ROM4[1222]<=26'd23462712;
ROM1[1223]<=26'd1944111; ROM2[1223]<=26'd11283136; ROM3[1223]<=26'd9755739; ROM4[1223]<=26'd23463993;
ROM1[1224]<=26'd1963117; ROM2[1224]<=26'd11291990; ROM3[1224]<=26'd9757992; ROM4[1224]<=26'd23470307;
ROM1[1225]<=26'd1977771; ROM2[1225]<=26'd11299304; ROM3[1225]<=26'd9757070; ROM4[1225]<=26'd23473680;
ROM1[1226]<=26'd1970102; ROM2[1226]<=26'd11294868; ROM3[1226]<=26'd9752805; ROM4[1226]<=26'd23469355;
ROM1[1227]<=26'd1958234; ROM2[1227]<=26'd11289134; ROM3[1227]<=26'd9750194; ROM4[1227]<=26'd23464725;
ROM1[1228]<=26'd1953501; ROM2[1228]<=26'd11292166; ROM3[1228]<=26'd9753362; ROM4[1228]<=26'd23465130;
ROM1[1229]<=26'd1956359; ROM2[1229]<=26'd11299765; ROM3[1229]<=26'd9763492; ROM4[1229]<=26'd23471715;
ROM1[1230]<=26'd1957187; ROM2[1230]<=26'd11303460; ROM3[1230]<=26'd9769574; ROM4[1230]<=26'd23475623;
ROM1[1231]<=26'd1952693; ROM2[1231]<=26'd11296421; ROM3[1231]<=26'd9762816; ROM4[1231]<=26'd23468056;
ROM1[1232]<=26'd1962464; ROM2[1232]<=26'd11294867; ROM3[1232]<=26'd9757474; ROM4[1232]<=26'd23467094;
ROM1[1233]<=26'd1973566; ROM2[1233]<=26'd11296517; ROM3[1233]<=26'd9752673; ROM4[1233]<=26'd23467785;
ROM1[1234]<=26'd1969036; ROM2[1234]<=26'd11291603; ROM3[1234]<=26'd9749293; ROM4[1234]<=26'd23464581;
ROM1[1235]<=26'd1965634; ROM2[1235]<=26'd11292278; ROM3[1235]<=26'd9754711; ROM4[1235]<=26'd23467309;
ROM1[1236]<=26'd1962642; ROM2[1236]<=26'd11295947; ROM3[1236]<=26'd9762926; ROM4[1236]<=26'd23471166;
ROM1[1237]<=26'd1955882; ROM2[1237]<=26'd11294453; ROM3[1237]<=26'd9764477; ROM4[1237]<=26'd23470060;
ROM1[1238]<=26'd1949295; ROM2[1238]<=26'd11293382; ROM3[1238]<=26'd9766588; ROM4[1238]<=26'd23469978;
ROM1[1239]<=26'd1950381; ROM2[1239]<=26'd11293530; ROM3[1239]<=26'd9766541; ROM4[1239]<=26'd23469624;
ROM1[1240]<=26'd1956737; ROM2[1240]<=26'd11290835; ROM3[1240]<=26'd9762227; ROM4[1240]<=26'd23467259;
ROM1[1241]<=26'd1970425; ROM2[1241]<=26'd11292355; ROM3[1241]<=26'd9757765; ROM4[1241]<=26'd23468517;
ROM1[1242]<=26'd1976343; ROM2[1242]<=26'd11293268; ROM3[1242]<=26'd9755513; ROM4[1242]<=26'd23468237;
ROM1[1243]<=26'd1972052; ROM2[1243]<=26'd11293231; ROM3[1243]<=26'd9758701; ROM4[1243]<=26'd23469403;
ROM1[1244]<=26'd1968276; ROM2[1244]<=26'd11294189; ROM3[1244]<=26'd9764666; ROM4[1244]<=26'd23472355;
ROM1[1245]<=26'd1964862; ROM2[1245]<=26'd11295027; ROM3[1245]<=26'd9768654; ROM4[1245]<=26'd23473427;
ROM1[1246]<=26'd1961173; ROM2[1246]<=26'd11298296; ROM3[1246]<=26'd9773143; ROM4[1246]<=26'd23476427;
ROM1[1247]<=26'd1962935; ROM2[1247]<=26'd11300215; ROM3[1247]<=26'd9775777; ROM4[1247]<=26'd23478836;
ROM1[1248]<=26'd1966337; ROM2[1248]<=26'd11299079; ROM3[1248]<=26'd9772478; ROM4[1248]<=26'd23476170;
ROM1[1249]<=26'd1969482; ROM2[1249]<=26'd11293503; ROM3[1249]<=26'd9761432; ROM4[1249]<=26'd23467740;
ROM1[1250]<=26'd1985724; ROM2[1250]<=26'd11301707; ROM3[1250]<=26'd9763065; ROM4[1250]<=26'd23473651;
ROM1[1251]<=26'd1994484; ROM2[1251]<=26'd11314890; ROM3[1251]<=26'd9773859; ROM4[1251]<=26'd23484206;
ROM1[1252]<=26'd1975209; ROM2[1252]<=26'd11303136; ROM3[1252]<=26'd9763795; ROM4[1252]<=26'd23472407;
ROM1[1253]<=26'd1958768; ROM2[1253]<=26'd11291759; ROM3[1253]<=26'd9758492; ROM4[1253]<=26'd23464302;
ROM1[1254]<=26'd1947899; ROM2[1254]<=26'd11285339; ROM3[1254]<=26'd9756217; ROM4[1254]<=26'd23461925;
ROM1[1255]<=26'd1937280; ROM2[1255]<=26'd11279956; ROM3[1255]<=26'd9750026; ROM4[1255]<=26'd23454944;
ROM1[1256]<=26'd1947540; ROM2[1256]<=26'd11288917; ROM3[1256]<=26'd9756676; ROM4[1256]<=26'd23462430;
ROM1[1257]<=26'd1965335; ROM2[1257]<=26'd11296647; ROM3[1257]<=26'd9759303; ROM4[1257]<=26'd23469579;
ROM1[1258]<=26'd1974957; ROM2[1258]<=26'd11296408; ROM3[1258]<=26'd9755229; ROM4[1258]<=26'd23467851;
ROM1[1259]<=26'd1972783; ROM2[1259]<=26'd11291804; ROM3[1259]<=26'd9753927; ROM4[1259]<=26'd23466938;
ROM1[1260]<=26'd1966961; ROM2[1260]<=26'd11292372; ROM3[1260]<=26'd9756456; ROM4[1260]<=26'd23467019;
ROM1[1261]<=26'd1960852; ROM2[1261]<=26'd11293141; ROM3[1261]<=26'd9758004; ROM4[1261]<=26'd23466565;
ROM1[1262]<=26'd1950027; ROM2[1262]<=26'd11286246; ROM3[1262]<=26'd9755410; ROM4[1262]<=26'd23461851;
ROM1[1263]<=26'd1939780; ROM2[1263]<=26'd11281195; ROM3[1263]<=26'd9756149; ROM4[1263]<=26'd23458321;
ROM1[1264]<=26'd1937478; ROM2[1264]<=26'd11279432; ROM3[1264]<=26'd9755543; ROM4[1264]<=26'd23457733;
ROM1[1265]<=26'd1946151; ROM2[1265]<=26'd11282052; ROM3[1265]<=26'd9753380; ROM4[1265]<=26'd23457224;
ROM1[1266]<=26'd1961029; ROM2[1266]<=26'd11286934; ROM3[1266]<=26'd9750364; ROM4[1266]<=26'd23456768;
ROM1[1267]<=26'd1958508; ROM2[1267]<=26'd11283354; ROM3[1267]<=26'd9741103; ROM4[1267]<=26'd23451005;
ROM1[1268]<=26'd1945963; ROM2[1268]<=26'd11276557; ROM3[1268]<=26'd9734627; ROM4[1268]<=26'd23444371;
ROM1[1269]<=26'd1937496; ROM2[1269]<=26'd11273565; ROM3[1269]<=26'd9735637; ROM4[1269]<=26'd23443280;
ROM1[1270]<=26'd1932937; ROM2[1270]<=26'd11275424; ROM3[1270]<=26'd9739469; ROM4[1270]<=26'd23446130;
ROM1[1271]<=26'd1930046; ROM2[1271]<=26'd11279701; ROM3[1271]<=26'd9745381; ROM4[1271]<=26'd23449298;
ROM1[1272]<=26'd1930116; ROM2[1272]<=26'd11279747; ROM3[1272]<=26'd9746696; ROM4[1272]<=26'd23450730;
ROM1[1273]<=26'd1940211; ROM2[1273]<=26'd11283028; ROM3[1273]<=26'd9748571; ROM4[1273]<=26'd23453983;
ROM1[1274]<=26'd1956569; ROM2[1274]<=26'd11286313; ROM3[1274]<=26'd9746698; ROM4[1274]<=26'd23455452;
ROM1[1275]<=26'd1962679; ROM2[1275]<=26'd11284239; ROM3[1275]<=26'd9740645; ROM4[1275]<=26'd23454349;
ROM1[1276]<=26'd1964130; ROM2[1276]<=26'd11289774; ROM3[1276]<=26'd9747899; ROM4[1276]<=26'd23459699;
ROM1[1277]<=26'd1959638; ROM2[1277]<=26'd11293609; ROM3[1277]<=26'd9756539; ROM4[1277]<=26'd23465056;
ROM1[1278]<=26'd1950340; ROM2[1278]<=26'd11289633; ROM3[1278]<=26'd9758559; ROM4[1278]<=26'd23463872;
ROM1[1279]<=26'd1946943; ROM2[1279]<=26'd11290109; ROM3[1279]<=26'd9762862; ROM4[1279]<=26'd23465669;
ROM1[1280]<=26'd1944538; ROM2[1280]<=26'd11290554; ROM3[1280]<=26'd9764534; ROM4[1280]<=26'd23465826;
ROM1[1281]<=26'd1948722; ROM2[1281]<=26'd11290738; ROM3[1281]<=26'd9764097; ROM4[1281]<=26'd23465856;
ROM1[1282]<=26'd1959947; ROM2[1282]<=26'd11293215; ROM3[1282]<=26'd9760054; ROM4[1282]<=26'd23466746;
ROM1[1283]<=26'd1973871; ROM2[1283]<=26'd11295840; ROM3[1283]<=26'd9757656; ROM4[1283]<=26'd23469665;
ROM1[1284]<=26'd1975381; ROM2[1284]<=26'd11298651; ROM3[1284]<=26'd9760781; ROM4[1284]<=26'd23473033;
ROM1[1285]<=26'd1971082; ROM2[1285]<=26'd11299842; ROM3[1285]<=26'd9766267; ROM4[1285]<=26'd23475235;
ROM1[1286]<=26'd1967199; ROM2[1286]<=26'd11299156; ROM3[1286]<=26'd9771092; ROM4[1286]<=26'd23475642;
ROM1[1287]<=26'd1959951; ROM2[1287]<=26'd11297554; ROM3[1287]<=26'd9771456; ROM4[1287]<=26'd23474656;
ROM1[1288]<=26'd1955099; ROM2[1288]<=26'd11298937; ROM3[1288]<=26'd9774410; ROM4[1288]<=26'd23476251;
ROM1[1289]<=26'd1955861; ROM2[1289]<=26'd11299516; ROM3[1289]<=26'd9772570; ROM4[1289]<=26'd23476256;
ROM1[1290]<=26'd1959188; ROM2[1290]<=26'd11296217; ROM3[1290]<=26'd9764813; ROM4[1290]<=26'd23472009;
ROM1[1291]<=26'd1974191; ROM2[1291]<=26'd11297653; ROM3[1291]<=26'd9763316; ROM4[1291]<=26'd23473440;
ROM1[1292]<=26'd1984676; ROM2[1292]<=26'd11300187; ROM3[1292]<=26'd9764662; ROM4[1292]<=26'd23476439;
ROM1[1293]<=26'd1981980; ROM2[1293]<=26'd11303032; ROM3[1293]<=26'd9769045; ROM4[1293]<=26'd23478520;
ROM1[1294]<=26'd1972613; ROM2[1294]<=26'd11300276; ROM3[1294]<=26'd9771858; ROM4[1294]<=26'd23477228;
ROM1[1295]<=26'd1963764; ROM2[1295]<=26'd11297545; ROM3[1295]<=26'd9770963; ROM4[1295]<=26'd23473073;
ROM1[1296]<=26'd1960382; ROM2[1296]<=26'd11300360; ROM3[1296]<=26'd9776102; ROM4[1296]<=26'd23475153;
ROM1[1297]<=26'd1957045; ROM2[1297]<=26'd11298642; ROM3[1297]<=26'd9776448; ROM4[1297]<=26'd23473815;
ROM1[1298]<=26'd1962032; ROM2[1298]<=26'd11299292; ROM3[1298]<=26'd9771690; ROM4[1298]<=26'd23471808;
ROM1[1299]<=26'd1973421; ROM2[1299]<=26'd11297595; ROM3[1299]<=26'd9761962; ROM4[1299]<=26'd23468205;
ROM1[1300]<=26'd1972467; ROM2[1300]<=26'd11289140; ROM3[1300]<=26'd9749291; ROM4[1300]<=26'd23460824;
ROM1[1301]<=26'd1967400; ROM2[1301]<=26'd11285388; ROM3[1301]<=26'd9747108; ROM4[1301]<=26'd23459320;
ROM1[1302]<=26'd1961897; ROM2[1302]<=26'd11286744; ROM3[1302]<=26'd9752077; ROM4[1302]<=26'd23461591;
ROM1[1303]<=26'd1958522; ROM2[1303]<=26'd11290780; ROM3[1303]<=26'd9758602; ROM4[1303]<=26'd23464381;
ROM1[1304]<=26'd1958558; ROM2[1304]<=26'd11295183; ROM3[1304]<=26'd9764522; ROM4[1304]<=26'd23468391;
ROM1[1305]<=26'd1957455; ROM2[1305]<=26'd11296230; ROM3[1305]<=26'd9766711; ROM4[1305]<=26'd23469277;
ROM1[1306]<=26'd1958181; ROM2[1306]<=26'd11293038; ROM3[1306]<=26'd9762054; ROM4[1306]<=26'd23466095;
ROM1[1307]<=26'd1965586; ROM2[1307]<=26'd11291486; ROM3[1307]<=26'd9755960; ROM4[1307]<=26'd23464371;
ROM1[1308]<=26'd1975707; ROM2[1308]<=26'd11291998; ROM3[1308]<=26'd9749561; ROM4[1308]<=26'd23462390;
ROM1[1309]<=26'd1971230; ROM2[1309]<=26'd11290133; ROM3[1309]<=26'd9745899; ROM4[1309]<=26'd23460810;
ROM1[1310]<=26'd1969034; ROM2[1310]<=26'd11294201; ROM3[1310]<=26'd9753365; ROM4[1310]<=26'd23466081;
ROM1[1311]<=26'd1969234; ROM2[1311]<=26'd11299491; ROM3[1311]<=26'd9762547; ROM4[1311]<=26'd23471056;
ROM1[1312]<=26'd1967219; ROM2[1312]<=26'd11303106; ROM3[1312]<=26'd9769729; ROM4[1312]<=26'd23476112;
ROM1[1313]<=26'd1966111; ROM2[1313]<=26'd11306151; ROM3[1313]<=26'd9774893; ROM4[1313]<=26'd23479778;
ROM1[1314]<=26'd1968545; ROM2[1314]<=26'd11309755; ROM3[1314]<=26'd9777520; ROM4[1314]<=26'd23481690;
ROM1[1315]<=26'd1970478; ROM2[1315]<=26'd11304829; ROM3[1315]<=26'd9767543; ROM4[1315]<=26'd23474967;
ROM1[1316]<=26'd1970293; ROM2[1316]<=26'd11292031; ROM3[1316]<=26'd9748714; ROM4[1316]<=26'd23461955;
ROM1[1317]<=26'd1972013; ROM2[1317]<=26'd11290133; ROM3[1317]<=26'd9745528; ROM4[1317]<=26'd23460825;
ROM1[1318]<=26'd1968970; ROM2[1318]<=26'd11290345; ROM3[1318]<=26'd9747101; ROM4[1318]<=26'd23460597;
ROM1[1319]<=26'd1965685; ROM2[1319]<=26'd11292937; ROM3[1319]<=26'd9751869; ROM4[1319]<=26'd23463448;
ROM1[1320]<=26'd1966850; ROM2[1320]<=26'd11299556; ROM3[1320]<=26'd9762526; ROM4[1320]<=26'd23470341;
ROM1[1321]<=26'd1956890; ROM2[1321]<=26'd11295453; ROM3[1321]<=26'd9763201; ROM4[1321]<=26'd23467404;
ROM1[1322]<=26'd1950592; ROM2[1322]<=26'd11291308; ROM3[1322]<=26'd9759089; ROM4[1322]<=26'd23465800;
ROM1[1323]<=26'd1956427; ROM2[1323]<=26'd11293001; ROM3[1323]<=26'd9758821; ROM4[1323]<=26'd23467251;
ROM1[1324]<=26'd1972586; ROM2[1324]<=26'd11297939; ROM3[1324]<=26'd9756707; ROM4[1324]<=26'd23469622;
ROM1[1325]<=26'd1987128; ROM2[1325]<=26'd11304829; ROM3[1325]<=26'd9757235; ROM4[1325]<=26'd23474943;
ROM1[1326]<=26'd1987662; ROM2[1326]<=26'd11306267; ROM3[1326]<=26'd9761166; ROM4[1326]<=26'd23477891;
ROM1[1327]<=26'd1978786; ROM2[1327]<=26'd11304262; ROM3[1327]<=26'd9764196; ROM4[1327]<=26'd23477600;
ROM1[1328]<=26'd1969219; ROM2[1328]<=26'd11300679; ROM3[1328]<=26'd9763831; ROM4[1328]<=26'd23474362;
ROM1[1329]<=26'd1961026; ROM2[1329]<=26'd11298315; ROM3[1329]<=26'd9764705; ROM4[1329]<=26'd23471728;
ROM1[1330]<=26'd1958216; ROM2[1330]<=26'd11299543; ROM3[1330]<=26'd9767148; ROM4[1330]<=26'd23471713;
ROM1[1331]<=26'd1963015; ROM2[1331]<=26'd11299752; ROM3[1331]<=26'd9766995; ROM4[1331]<=26'd23470499;
ROM1[1332]<=26'd1973955; ROM2[1332]<=26'd11298874; ROM3[1332]<=26'd9764567; ROM4[1332]<=26'd23471016;
ROM1[1333]<=26'd1982920; ROM2[1333]<=26'd11297853; ROM3[1333]<=26'd9760236; ROM4[1333]<=26'd23470235;
ROM1[1334]<=26'd1979820; ROM2[1334]<=26'd11295451; ROM3[1334]<=26'd9761500; ROM4[1334]<=26'd23469081;
ROM1[1335]<=26'd1973909; ROM2[1335]<=26'd11294876; ROM3[1335]<=26'd9765677; ROM4[1335]<=26'd23469659;
ROM1[1336]<=26'd1966121; ROM2[1336]<=26'd11293348; ROM3[1336]<=26'd9767646; ROM4[1336]<=26'd23467349;
ROM1[1337]<=26'd1958083; ROM2[1337]<=26'd11289479; ROM3[1337]<=26'd9766108; ROM4[1337]<=26'd23463503;
ROM1[1338]<=26'd1951804; ROM2[1338]<=26'd11288684; ROM3[1338]<=26'd9766554; ROM4[1338]<=26'd23463200;
ROM1[1339]<=26'd1950745; ROM2[1339]<=26'd11289412; ROM3[1339]<=26'd9763880; ROM4[1339]<=26'd23464389;
ROM1[1340]<=26'd1959151; ROM2[1340]<=26'd11291599; ROM3[1340]<=26'd9761391; ROM4[1340]<=26'd23464618;
ROM1[1341]<=26'd1981835; ROM2[1341]<=26'd11303392; ROM3[1341]<=26'd9765011; ROM4[1341]<=26'd23472629;
ROM1[1342]<=26'd1985363; ROM2[1342]<=26'd11303335; ROM3[1342]<=26'd9762162; ROM4[1342]<=26'd23472919;
ROM1[1343]<=26'd1975347; ROM2[1343]<=26'd11298180; ROM3[1343]<=26'd9761056; ROM4[1343]<=26'd23469696;
ROM1[1344]<=26'd1965818; ROM2[1344]<=26'd11296360; ROM3[1344]<=26'd9761750; ROM4[1344]<=26'd23468504;
ROM1[1345]<=26'd1953158; ROM2[1345]<=26'd11287360; ROM3[1345]<=26'd9756221; ROM4[1345]<=26'd23460286;
ROM1[1346]<=26'd1953923; ROM2[1346]<=26'd11293985; ROM3[1346]<=26'd9763945; ROM4[1346]<=26'd23466518;
ROM1[1347]<=26'd1953490; ROM2[1347]<=26'd11295303; ROM3[1347]<=26'd9765102; ROM4[1347]<=26'd23467263;
ROM1[1348]<=26'd1956318; ROM2[1348]<=26'd11294097; ROM3[1348]<=26'd9761324; ROM4[1348]<=26'd23464134;
ROM1[1349]<=26'd1970098; ROM2[1349]<=26'd11297314; ROM3[1349]<=26'd9758652; ROM4[1349]<=26'd23467300;
ROM1[1350]<=26'd1984381; ROM2[1350]<=26'd11302759; ROM3[1350]<=26'd9759315; ROM4[1350]<=26'd23471262;
ROM1[1351]<=26'd1985785; ROM2[1351]<=26'd11308814; ROM3[1351]<=26'd9764588; ROM4[1351]<=26'd23475509;
ROM1[1352]<=26'd1971813; ROM2[1352]<=26'd11301347; ROM3[1352]<=26'd9758984; ROM4[1352]<=26'd23468858;
ROM1[1353]<=26'd1962147; ROM2[1353]<=26'd11297973; ROM3[1353]<=26'd9757491; ROM4[1353]<=26'd23465999;
ROM1[1354]<=26'd1948804; ROM2[1354]<=26'd11292498; ROM3[1354]<=26'd9756110; ROM4[1354]<=26'd23462618;
ROM1[1355]<=26'd1941111; ROM2[1355]<=26'd11287115; ROM3[1355]<=26'd9753253; ROM4[1355]<=26'd23457488;
ROM1[1356]<=26'd1944960; ROM2[1356]<=26'd11288511; ROM3[1356]<=26'd9752577; ROM4[1356]<=26'd23458379;
ROM1[1357]<=26'd1953640; ROM2[1357]<=26'd11287100; ROM3[1357]<=26'd9746266; ROM4[1357]<=26'd23456213;
ROM1[1358]<=26'd1961364; ROM2[1358]<=26'd11283475; ROM3[1358]<=26'd9736231; ROM4[1358]<=26'd23449747;
ROM1[1359]<=26'd1959662; ROM2[1359]<=26'd11282952; ROM3[1359]<=26'd9736330; ROM4[1359]<=26'd23448569;
ROM1[1360]<=26'd1960042; ROM2[1360]<=26'd11288167; ROM3[1360]<=26'd9748159; ROM4[1360]<=26'd23456926;
ROM1[1361]<=26'd1955990; ROM2[1361]<=26'd11288697; ROM3[1361]<=26'd9754061; ROM4[1361]<=26'd23459879;
ROM1[1362]<=26'd1946474; ROM2[1362]<=26'd11284063; ROM3[1362]<=26'd9752380; ROM4[1362]<=26'd23456295;
ROM1[1363]<=26'd1942022; ROM2[1363]<=26'd11283397; ROM3[1363]<=26'd9755800; ROM4[1363]<=26'd23458181;
ROM1[1364]<=26'd1945973; ROM2[1364]<=26'd11287261; ROM3[1364]<=26'd9759529; ROM4[1364]<=26'd23461859;
ROM1[1365]<=26'd1960013; ROM2[1365]<=26'd11295766; ROM3[1365]<=26'd9764015; ROM4[1365]<=26'd23468248;
ROM1[1366]<=26'd1984782; ROM2[1366]<=26'd11307274; ROM3[1366]<=26'd9771886; ROM4[1366]<=26'd23480085;
ROM1[1367]<=26'd1990751; ROM2[1367]<=26'd11310059; ROM3[1367]<=26'd9773081; ROM4[1367]<=26'd23483787;
ROM1[1368]<=26'd1969247; ROM2[1368]<=26'd11294546; ROM3[1368]<=26'd9762314; ROM4[1368]<=26'd23470599;
ROM1[1369]<=26'd1953844; ROM2[1369]<=26'd11286004; ROM3[1369]<=26'd9760205; ROM4[1369]<=26'd23463422;
ROM1[1370]<=26'd1946413; ROM2[1370]<=26'd11284881; ROM3[1370]<=26'd9761422; ROM4[1370]<=26'd23462566;
ROM1[1371]<=26'd1945451; ROM2[1371]<=26'd11287867; ROM3[1371]<=26'd9765804; ROM4[1371]<=26'd23465674;
ROM1[1372]<=26'd1959913; ROM2[1372]<=26'd11301960; ROM3[1372]<=26'd9779589; ROM4[1372]<=26'd23478933;
ROM1[1373]<=26'd1973181; ROM2[1373]<=26'd11309151; ROM3[1373]<=26'd9784119; ROM4[1373]<=26'd23485099;
ROM1[1374]<=26'd1976308; ROM2[1374]<=26'd11300358; ROM3[1374]<=26'd9771682; ROM4[1374]<=26'd23474797;
ROM1[1375]<=26'd1976778; ROM2[1375]<=26'd11295124; ROM3[1375]<=26'd9762216; ROM4[1375]<=26'd23468880;
ROM1[1376]<=26'd1973604; ROM2[1376]<=26'd11293431; ROM3[1376]<=26'd9760975; ROM4[1376]<=26'd23469083;
ROM1[1377]<=26'd1966340; ROM2[1377]<=26'd11292064; ROM3[1377]<=26'd9762060; ROM4[1377]<=26'd23469019;
ROM1[1378]<=26'd1963869; ROM2[1378]<=26'd11295382; ROM3[1378]<=26'd9765810; ROM4[1378]<=26'd23472728;
ROM1[1379]<=26'd1959374; ROM2[1379]<=26'd11294617; ROM3[1379]<=26'd9769963; ROM4[1379]<=26'd23474446;
ROM1[1380]<=26'd1957555; ROM2[1380]<=26'd11297753; ROM3[1380]<=26'd9774130; ROM4[1380]<=26'd23476158;
ROM1[1381]<=26'd1961060; ROM2[1381]<=26'd11298999; ROM3[1381]<=26'd9772460; ROM4[1381]<=26'd23475470;
ROM1[1382]<=26'd1974957; ROM2[1382]<=26'd11304788; ROM3[1382]<=26'd9772342; ROM4[1382]<=26'd23479276;
ROM1[1383]<=26'd1990606; ROM2[1383]<=26'd11309308; ROM3[1383]<=26'd9770503; ROM4[1383]<=26'd23483838;
ROM1[1384]<=26'd1985954; ROM2[1384]<=26'd11304677; ROM3[1384]<=26'd9767963; ROM4[1384]<=26'd23480939;
ROM1[1385]<=26'd1975053; ROM2[1385]<=26'd11300532; ROM3[1385]<=26'd9769496; ROM4[1385]<=26'd23479214;
ROM1[1386]<=26'd1967652; ROM2[1386]<=26'd11296394; ROM3[1386]<=26'd9771570; ROM4[1386]<=26'd23477706;
ROM1[1387]<=26'd1961755; ROM2[1387]<=26'd11293984; ROM3[1387]<=26'd9774304; ROM4[1387]<=26'd23476167;
ROM1[1388]<=26'd1956901; ROM2[1388]<=26'd11293869; ROM3[1388]<=26'd9776766; ROM4[1388]<=26'd23477542;
ROM1[1389]<=26'd1956425; ROM2[1389]<=26'd11292493; ROM3[1389]<=26'd9774717; ROM4[1389]<=26'd23476214;
ROM1[1390]<=26'd1962585; ROM2[1390]<=26'd11292640; ROM3[1390]<=26'd9769976; ROM4[1390]<=26'd23473597;
ROM1[1391]<=26'd1973657; ROM2[1391]<=26'd11294006; ROM3[1391]<=26'd9763924; ROM4[1391]<=26'd23471977;
ROM1[1392]<=26'd1977954; ROM2[1392]<=26'd11294104; ROM3[1392]<=26'd9761553; ROM4[1392]<=26'd23471797;
ROM1[1393]<=26'd1973450; ROM2[1393]<=26'd11295241; ROM3[1393]<=26'd9764776; ROM4[1393]<=26'd23472810;
ROM1[1394]<=26'd1963182; ROM2[1394]<=26'd11293031; ROM3[1394]<=26'd9767486; ROM4[1394]<=26'd23471680;
ROM1[1395]<=26'd1955639; ROM2[1395]<=26'd11290864; ROM3[1395]<=26'd9767256; ROM4[1395]<=26'd23469512;
ROM1[1396]<=26'd1956848; ROM2[1396]<=26'd11299874; ROM3[1396]<=26'd9776982; ROM4[1396]<=26'd23477376;
ROM1[1397]<=26'd1966158; ROM2[1397]<=26'd11311523; ROM3[1397]<=26'd9786992; ROM4[1397]<=26'd23486603;
ROM1[1398]<=26'd1970420; ROM2[1398]<=26'd11310204; ROM3[1398]<=26'd9780031; ROM4[1398]<=26'd23482670;
ROM1[1399]<=26'd1964379; ROM2[1399]<=26'd11290645; ROM3[1399]<=26'd9755407; ROM4[1399]<=26'd23462429;
ROM1[1400]<=26'd1958897; ROM2[1400]<=26'd11275390; ROM3[1400]<=26'd9737646; ROM4[1400]<=26'd23446888;
ROM1[1401]<=26'd1950458; ROM2[1401]<=26'd11269570; ROM3[1401]<=26'd9735702; ROM4[1401]<=26'd23443699;
ROM1[1402]<=26'd1941088; ROM2[1402]<=26'd11268492; ROM3[1402]<=26'd9739279; ROM4[1402]<=26'd23444629;
ROM1[1403]<=26'd1942081; ROM2[1403]<=26'd11276521; ROM3[1403]<=26'd9750822; ROM4[1403]<=26'd23452389;
ROM1[1404]<=26'd1939193; ROM2[1404]<=26'd11279330; ROM3[1404]<=26'd9754605; ROM4[1404]<=26'd23454619;
ROM1[1405]<=26'd1933984; ROM2[1405]<=26'd11277347; ROM3[1405]<=26'd9752050; ROM4[1405]<=26'd23452328;
ROM1[1406]<=26'd1940928; ROM2[1406]<=26'd11281167; ROM3[1406]<=26'd9753613; ROM4[1406]<=26'd23454636;
ROM1[1407]<=26'd1957116; ROM2[1407]<=26'd11288823; ROM3[1407]<=26'd9754645; ROM4[1407]<=26'd23460117;
ROM1[1408]<=26'd1970407; ROM2[1408]<=26'd11291242; ROM3[1408]<=26'd9753562; ROM4[1408]<=26'd23463258;
ROM1[1409]<=26'd1970762; ROM2[1409]<=26'd11293009; ROM3[1409]<=26'd9754161; ROM4[1409]<=26'd23464979;
ROM1[1410]<=26'd1967727; ROM2[1410]<=26'd11295894; ROM3[1410]<=26'd9757667; ROM4[1410]<=26'd23467858;
ROM1[1411]<=26'd1958405; ROM2[1411]<=26'd11292353; ROM3[1411]<=26'd9758700; ROM4[1411]<=26'd23466706;
ROM1[1412]<=26'd1947823; ROM2[1412]<=26'd11287289; ROM3[1412]<=26'd9756702; ROM4[1412]<=26'd23462445;
ROM1[1413]<=26'd1944707; ROM2[1413]<=26'd11288496; ROM3[1413]<=26'd9759248; ROM4[1413]<=26'd23463271;
ROM1[1414]<=26'd1949045; ROM2[1414]<=26'd11290590; ROM3[1414]<=26'd9762669; ROM4[1414]<=26'd23466241;
ROM1[1415]<=26'd1962365; ROM2[1415]<=26'd11293715; ROM3[1415]<=26'd9764100; ROM4[1415]<=26'd23470540;
ROM1[1416]<=26'd1978322; ROM2[1416]<=26'd11297393; ROM3[1416]<=26'd9761548; ROM4[1416]<=26'd23473503;
ROM1[1417]<=26'd1975753; ROM2[1417]<=26'd11291676; ROM3[1417]<=26'd9753557; ROM4[1417]<=26'd23466140;
ROM1[1418]<=26'd1968499; ROM2[1418]<=26'd11289448; ROM3[1418]<=26'd9755111; ROM4[1418]<=26'd23464908;
ROM1[1419]<=26'd1969718; ROM2[1419]<=26'd11297226; ROM3[1419]<=26'd9767926; ROM4[1419]<=26'd23473100;
ROM1[1420]<=26'd1964518; ROM2[1420]<=26'd11298733; ROM3[1420]<=26'd9773575; ROM4[1420]<=26'd23475239;
ROM1[1421]<=26'd1955222; ROM2[1421]<=26'd11293763; ROM3[1421]<=26'd9774286; ROM4[1421]<=26'd23472724;
ROM1[1422]<=26'd1946662; ROM2[1422]<=26'd11287554; ROM3[1422]<=26'd9765851; ROM4[1422]<=26'd23465311;
ROM1[1423]<=26'd1947208; ROM2[1423]<=26'd11283059; ROM3[1423]<=26'd9756531; ROM4[1423]<=26'd23459108;
ROM1[1424]<=26'd1962975; ROM2[1424]<=26'd11285549; ROM3[1424]<=26'd9754447; ROM4[1424]<=26'd23458893;
ROM1[1425]<=26'd1970894; ROM2[1425]<=26'd11287153; ROM3[1425]<=26'd9752925; ROM4[1425]<=26'd23461608;
ROM1[1426]<=26'd1967715; ROM2[1426]<=26'd11287221; ROM3[1426]<=26'd9756555; ROM4[1426]<=26'd23464062;
ROM1[1427]<=26'd1962327; ROM2[1427]<=26'd11289881; ROM3[1427]<=26'd9761631; ROM4[1427]<=26'd23465651;
ROM1[1428]<=26'd1959589; ROM2[1428]<=26'd11292434; ROM3[1428]<=26'd9766423; ROM4[1428]<=26'd23469365;
ROM1[1429]<=26'd1957927; ROM2[1429]<=26'd11292996; ROM3[1429]<=26'd9772193; ROM4[1429]<=26'd23472519;
ROM1[1430]<=26'd1956906; ROM2[1430]<=26'd11293739; ROM3[1430]<=26'd9776083; ROM4[1430]<=26'd23474000;
ROM1[1431]<=26'd1959389; ROM2[1431]<=26'd11293599; ROM3[1431]<=26'd9773895; ROM4[1431]<=26'd23472885;
ROM1[1432]<=26'd1967724; ROM2[1432]<=26'd11292484; ROM3[1432]<=26'd9766520; ROM4[1432]<=26'd23471193;
ROM1[1433]<=26'd1978679; ROM2[1433]<=26'd11295152; ROM3[1433]<=26'd9762432; ROM4[1433]<=26'd23471923;
ROM1[1434]<=26'd1978953; ROM2[1434]<=26'd11297489; ROM3[1434]<=26'd9764326; ROM4[1434]<=26'd23474024;
ROM1[1435]<=26'd1973374; ROM2[1435]<=26'd11297785; ROM3[1435]<=26'd9768706; ROM4[1435]<=26'd23476504;
ROM1[1436]<=26'd1963960; ROM2[1436]<=26'd11295294; ROM3[1436]<=26'd9770011; ROM4[1436]<=26'd23474567;
ROM1[1437]<=26'd1954362; ROM2[1437]<=26'd11291173; ROM3[1437]<=26'd9769352; ROM4[1437]<=26'd23471341;
ROM1[1438]<=26'd1949575; ROM2[1438]<=26'd11292167; ROM3[1438]<=26'd9770535; ROM4[1438]<=26'd23471821;
ROM1[1439]<=26'd1952052; ROM2[1439]<=26'd11295502; ROM3[1439]<=26'd9772837; ROM4[1439]<=26'd23474161;
ROM1[1440]<=26'd1961047; ROM2[1440]<=26'd11296749; ROM3[1440]<=26'd9768248; ROM4[1440]<=26'd23473335;
ROM1[1441]<=26'd1980718; ROM2[1441]<=26'd11305202; ROM3[1441]<=26'd9766237; ROM4[1441]<=26'd23476417;
ROM1[1442]<=26'd1986370; ROM2[1442]<=26'd11307596; ROM3[1442]<=26'd9768804; ROM4[1442]<=26'd23479919;
ROM1[1443]<=26'd1974285; ROM2[1443]<=26'd11302375; ROM3[1443]<=26'd9765288; ROM4[1443]<=26'd23476006;
ROM1[1444]<=26'd1960021; ROM2[1444]<=26'd11294969; ROM3[1444]<=26'd9761132; ROM4[1444]<=26'd23468410;
ROM1[1445]<=26'd1952530; ROM2[1445]<=26'd11290551; ROM3[1445]<=26'd9762353; ROM4[1445]<=26'd23467152;
ROM1[1446]<=26'd1943752; ROM2[1446]<=26'd11285969; ROM3[1446]<=26'd9761136; ROM4[1446]<=26'd23463800;
ROM1[1447]<=26'd1942988; ROM2[1447]<=26'd11285624; ROM3[1447]<=26'd9760101; ROM4[1447]<=26'd23462798;
ROM1[1448]<=26'd1952737; ROM2[1448]<=26'd11290452; ROM3[1448]<=26'd9760617; ROM4[1448]<=26'd23466275;
ROM1[1449]<=26'd1961291; ROM2[1449]<=26'd11288836; ROM3[1449]<=26'd9751361; ROM4[1449]<=26'd23462757;
ROM1[1450]<=26'd1965593; ROM2[1450]<=26'd11285243; ROM3[1450]<=26'd9741936; ROM4[1450]<=26'd23456657;
ROM1[1451]<=26'd1957356; ROM2[1451]<=26'd11279419; ROM3[1451]<=26'd9737916; ROM4[1451]<=26'd23451136;
ROM1[1452]<=26'd1948168; ROM2[1452]<=26'd11278138; ROM3[1452]<=26'd9742402; ROM4[1452]<=26'd23451786;
ROM1[1453]<=26'd1943916; ROM2[1453]<=26'd11279622; ROM3[1453]<=26'd9747368; ROM4[1453]<=26'd23453837;
ROM1[1454]<=26'd1931567; ROM2[1454]<=26'd11274548; ROM3[1454]<=26'd9744708; ROM4[1454]<=26'd23449158;
ROM1[1455]<=26'd1927661; ROM2[1455]<=26'd11273550; ROM3[1455]<=26'd9746255; ROM4[1455]<=26'd23449371;
ROM1[1456]<=26'd1933794; ROM2[1456]<=26'd11277520; ROM3[1456]<=26'd9749088; ROM4[1456]<=26'd23452984;
ROM1[1457]<=26'd1942905; ROM2[1457]<=26'd11277083; ROM3[1457]<=26'd9744767; ROM4[1457]<=26'd23450862;
ROM1[1458]<=26'd1955150; ROM2[1458]<=26'd11279412; ROM3[1458]<=26'd9742956; ROM4[1458]<=26'd23453944;
ROM1[1459]<=26'd1955230; ROM2[1459]<=26'd11281967; ROM3[1459]<=26'd9744549; ROM4[1459]<=26'd23456046;
ROM1[1460]<=26'd1948096; ROM2[1460]<=26'd11281643; ROM3[1460]<=26'd9748004; ROM4[1460]<=26'd23456619;
ROM1[1461]<=26'd1942308; ROM2[1461]<=26'd11281728; ROM3[1461]<=26'd9753545; ROM4[1461]<=26'd23458379;
ROM1[1462]<=26'd1943215; ROM2[1462]<=26'd11285257; ROM3[1462]<=26'd9761299; ROM4[1462]<=26'd23462237;
ROM1[1463]<=26'd1942635; ROM2[1463]<=26'd11288971; ROM3[1463]<=26'd9768141; ROM4[1463]<=26'd23468190;
ROM1[1464]<=26'd1951863; ROM2[1464]<=26'd11297075; ROM3[1464]<=26'd9775759; ROM4[1464]<=26'd23476231;
ROM1[1465]<=26'd1960960; ROM2[1465]<=26'd11297870; ROM3[1465]<=26'd9771996; ROM4[1465]<=26'd23474472;
ROM1[1466]<=26'd1965666; ROM2[1466]<=26'd11290160; ROM3[1466]<=26'd9759407; ROM4[1466]<=26'd23466070;
ROM1[1467]<=26'd1975177; ROM2[1467]<=26'd11295252; ROM3[1467]<=26'd9765066; ROM4[1467]<=26'd23471179;
ROM1[1468]<=26'd1975637; ROM2[1468]<=26'd11300359; ROM3[1468]<=26'd9773835; ROM4[1468]<=26'd23477832;
ROM1[1469]<=26'd1971597; ROM2[1469]<=26'd11301396; ROM3[1469]<=26'd9780525; ROM4[1469]<=26'd23481763;
ROM1[1470]<=26'd1965277; ROM2[1470]<=26'd11299488; ROM3[1470]<=26'd9781277; ROM4[1470]<=26'd23480127;
ROM1[1471]<=26'd1949568; ROM2[1471]<=26'd11289351; ROM3[1471]<=26'd9774674; ROM4[1471]<=26'd23470693;
ROM1[1472]<=26'd1936781; ROM2[1472]<=26'd11277740; ROM3[1472]<=26'd9763346; ROM4[1472]<=26'd23459467;
ROM1[1473]<=26'd1939510; ROM2[1473]<=26'd11274895; ROM3[1473]<=26'd9756741; ROM4[1473]<=26'd23456227;
ROM1[1474]<=26'd1956520; ROM2[1474]<=26'd11280575; ROM3[1474]<=26'd9757240; ROM4[1474]<=26'd23459810;
ROM1[1475]<=26'd1967483; ROM2[1475]<=26'd11285364; ROM3[1475]<=26'd9756582; ROM4[1475]<=26'd23462872;
ROM1[1476]<=26'd1966888; ROM2[1476]<=26'd11287677; ROM3[1476]<=26'd9760729; ROM4[1476]<=26'd23465202;
ROM1[1477]<=26'd1962166; ROM2[1477]<=26'd11290291; ROM3[1477]<=26'd9768231; ROM4[1477]<=26'd23469009;
ROM1[1478]<=26'd1959926; ROM2[1478]<=26'd11294390; ROM3[1478]<=26'd9775713; ROM4[1478]<=26'd23474876;
ROM1[1479]<=26'd1953315; ROM2[1479]<=26'd11291343; ROM3[1479]<=26'd9776184; ROM4[1479]<=26'd23473909;
ROM1[1480]<=26'd1946666; ROM2[1480]<=26'd11285663; ROM3[1480]<=26'd9772827; ROM4[1480]<=26'd23469669;
ROM1[1481]<=26'd1945157; ROM2[1481]<=26'd11283285; ROM3[1481]<=26'd9767384; ROM4[1481]<=26'd23466442;
ROM1[1482]<=26'd1953050; ROM2[1482]<=26'd11283770; ROM3[1482]<=26'd9760849; ROM4[1482]<=26'd23465997;
ROM1[1483]<=26'd1964116; ROM2[1483]<=26'd11284872; ROM3[1483]<=26'd9755380; ROM4[1483]<=26'd23464992;
ROM1[1484]<=26'd1962325; ROM2[1484]<=26'd11284871; ROM3[1484]<=26'd9754897; ROM4[1484]<=26'd23464161;
ROM1[1485]<=26'd1956765; ROM2[1485]<=26'd11286109; ROM3[1485]<=26'd9759547; ROM4[1485]<=26'd23467322;
ROM1[1486]<=26'd1954494; ROM2[1486]<=26'd11288889; ROM3[1486]<=26'd9766475; ROM4[1486]<=26'd23471741;
ROM1[1487]<=26'd1951647; ROM2[1487]<=26'd11290781; ROM3[1487]<=26'd9772548; ROM4[1487]<=26'd23475638;
ROM1[1488]<=26'd1944884; ROM2[1488]<=26'd11290278; ROM3[1488]<=26'd9774940; ROM4[1488]<=26'd23476848;
ROM1[1489]<=26'd1939935; ROM2[1489]<=26'd11284989; ROM3[1489]<=26'd9770328; ROM4[1489]<=26'd23469766;
ROM1[1490]<=26'd1947949; ROM2[1490]<=26'd11285063; ROM3[1490]<=26'd9767100; ROM4[1490]<=26'd23467105;
ROM1[1491]<=26'd1966711; ROM2[1491]<=26'd11294245; ROM3[1491]<=26'd9769932; ROM4[1491]<=26'd23474920;
ROM1[1492]<=26'd1969631; ROM2[1492]<=26'd11294447; ROM3[1492]<=26'd9768445; ROM4[1492]<=26'd23475510;
ROM1[1493]<=26'd1956693; ROM2[1493]<=26'd11286539; ROM3[1493]<=26'd9762070; ROM4[1493]<=26'd23467704;
ROM1[1494]<=26'd1946120; ROM2[1494]<=26'd11283745; ROM3[1494]<=26'd9760433; ROM4[1494]<=26'd23464707;
ROM1[1495]<=26'd1941700; ROM2[1495]<=26'd11282903; ROM3[1495]<=26'd9762519; ROM4[1495]<=26'd23463753;
ROM1[1496]<=26'd1937265; ROM2[1496]<=26'd11282488; ROM3[1496]<=26'd9765090; ROM4[1496]<=26'd23464391;
ROM1[1497]<=26'd1935507; ROM2[1497]<=26'd11282286; ROM3[1497]<=26'd9764989; ROM4[1497]<=26'd23464165;
ROM1[1498]<=26'd1937981; ROM2[1498]<=26'd11279510; ROM3[1498]<=26'd9760160; ROM4[1498]<=26'd23460270;
ROM1[1499]<=26'd1946673; ROM2[1499]<=26'd11277949; ROM3[1499]<=26'd9751423; ROM4[1499]<=26'd23456301;
ROM1[1500]<=26'd1953746; ROM2[1500]<=26'd11280471; ROM3[1500]<=26'd9746806; ROM4[1500]<=26'd23454419;
ROM1[1501]<=26'd1955660; ROM2[1501]<=26'd11285202; ROM3[1501]<=26'd9751966; ROM4[1501]<=26'd23459520;
ROM1[1502]<=26'd1951223; ROM2[1502]<=26'd11284352; ROM3[1502]<=26'd9756213; ROM4[1502]<=26'd23462543;
ROM1[1503]<=26'd1944262; ROM2[1503]<=26'd11282705; ROM3[1503]<=26'd9758634; ROM4[1503]<=26'd23463261;
ROM1[1504]<=26'd1940558; ROM2[1504]<=26'd11283629; ROM3[1504]<=26'd9762666; ROM4[1504]<=26'd23466098;
ROM1[1505]<=26'd1941105; ROM2[1505]<=26'd11286798; ROM3[1505]<=26'd9766066; ROM4[1505]<=26'd23467936;
ROM1[1506]<=26'd1940981; ROM2[1506]<=26'd11284056; ROM3[1506]<=26'd9761072; ROM4[1506]<=26'd23462333;
ROM1[1507]<=26'd1947098; ROM2[1507]<=26'd11279110; ROM3[1507]<=26'd9750698; ROM4[1507]<=26'd23455248;
ROM1[1508]<=26'd1956566; ROM2[1508]<=26'd11276469; ROM3[1508]<=26'd9746151; ROM4[1508]<=26'd23453352;
ROM1[1509]<=26'd1954182; ROM2[1509]<=26'd11276027; ROM3[1509]<=26'd9747613; ROM4[1509]<=26'd23454720;
ROM1[1510]<=26'd1948629; ROM2[1510]<=26'd11278005; ROM3[1510]<=26'd9752505; ROM4[1510]<=26'd23457317;
ROM1[1511]<=26'd1946997; ROM2[1511]<=26'd11282664; ROM3[1511]<=26'd9761523; ROM4[1511]<=26'd23462680;
ROM1[1512]<=26'd1953307; ROM2[1512]<=26'd11293278; ROM3[1512]<=26'd9774209; ROM4[1512]<=26'd23473008;
ROM1[1513]<=26'd1958751; ROM2[1513]<=26'd11301854; ROM3[1513]<=26'd9786121; ROM4[1513]<=26'd23481443;
ROM1[1514]<=26'd1953524; ROM2[1514]<=26'd11297060; ROM3[1514]<=26'd9780473; ROM4[1514]<=26'd23476199;
ROM1[1515]<=26'd1948871; ROM2[1515]<=26'd11283720; ROM3[1515]<=26'd9762227; ROM4[1515]<=26'd23462019;
ROM1[1516]<=26'd1955692; ROM2[1516]<=26'd11278197; ROM3[1516]<=26'd9751319; ROM4[1516]<=26'd23455603;
ROM1[1517]<=26'd1952182; ROM2[1517]<=26'd11272055; ROM3[1517]<=26'd9741133; ROM4[1517]<=26'd23450775;
ROM1[1518]<=26'd1948811; ROM2[1518]<=26'd11272815; ROM3[1518]<=26'd9745279; ROM4[1518]<=26'd23453050;
ROM1[1519]<=26'd1949540; ROM2[1519]<=26'd11282519; ROM3[1519]<=26'd9760258; ROM4[1519]<=26'd23464400;
ROM1[1520]<=26'd1939655; ROM2[1520]<=26'd11279630; ROM3[1520]<=26'd9758401; ROM4[1520]<=26'd23462009;
ROM1[1521]<=26'd1925684; ROM2[1521]<=26'd11270266; ROM3[1521]<=26'd9752158; ROM4[1521]<=26'd23452773;
ROM1[1522]<=26'd1922972; ROM2[1522]<=26'd11270290; ROM3[1522]<=26'd9753126; ROM4[1522]<=26'd23453008;
ROM1[1523]<=26'd1926578; ROM2[1523]<=26'd11268305; ROM3[1523]<=26'd9744413; ROM4[1523]<=26'd23447941;
ROM1[1524]<=26'd1933509; ROM2[1524]<=26'd11261901; ROM3[1524]<=26'd9731221; ROM4[1524]<=26'd23439202;
ROM1[1525]<=26'd1942575; ROM2[1525]<=26'd11264024; ROM3[1525]<=26'd9730219; ROM4[1525]<=26'd23441253;
ROM1[1526]<=26'd1947592; ROM2[1526]<=26'd11272050; ROM3[1526]<=26'd9739730; ROM4[1526]<=26'd23451366;
ROM1[1527]<=26'd1952590; ROM2[1527]<=26'd11281277; ROM3[1527]<=26'd9755318; ROM4[1527]<=26'd23462141;
ROM1[1528]<=26'd1960422; ROM2[1528]<=26'd11293580; ROM3[1528]<=26'd9770275; ROM4[1528]<=26'd23474740;
ROM1[1529]<=26'd1958529; ROM2[1529]<=26'd11298062; ROM3[1529]<=26'd9775614; ROM4[1529]<=26'd23478854;
ROM1[1530]<=26'd1951640; ROM2[1530]<=26'd11296168; ROM3[1530]<=26'd9774431; ROM4[1530]<=26'd23474994;
ROM1[1531]<=26'd1951596; ROM2[1531]<=26'd11295198; ROM3[1531]<=26'd9772647; ROM4[1531]<=26'd23474894;
ROM1[1532]<=26'd1967422; ROM2[1532]<=26'd11301421; ROM3[1532]<=26'd9777172; ROM4[1532]<=26'd23480798;
ROM1[1533]<=26'd1984314; ROM2[1533]<=26'd11307129; ROM3[1533]<=26'd9780630; ROM4[1533]<=26'd23484701;
ROM1[1534]<=26'd1977286; ROM2[1534]<=26'd11298869; ROM3[1534]<=26'd9773480; ROM4[1534]<=26'd23477826;
ROM1[1535]<=26'd1965688; ROM2[1535]<=26'd11291904; ROM3[1535]<=26'd9770793; ROM4[1535]<=26'd23472314;
ROM1[1536]<=26'd1958076; ROM2[1536]<=26'd11291056; ROM3[1536]<=26'd9774187; ROM4[1536]<=26'd23472152;
ROM1[1537]<=26'd1951578; ROM2[1537]<=26'd11289728; ROM3[1537]<=26'd9776591; ROM4[1537]<=26'd23472798;
ROM1[1538]<=26'd1945312; ROM2[1538]<=26'd11290060; ROM3[1538]<=26'd9778772; ROM4[1538]<=26'd23474839;
ROM1[1539]<=26'd1946634; ROM2[1539]<=26'd11291589; ROM3[1539]<=26'd9780995; ROM4[1539]<=26'd23476771;
ROM1[1540]<=26'd1955613; ROM2[1540]<=26'd11291882; ROM3[1540]<=26'd9777126; ROM4[1540]<=26'd23476127;
ROM1[1541]<=26'd1966541; ROM2[1541]<=26'd11290939; ROM3[1541]<=26'd9767679; ROM4[1541]<=26'd23473417;
ROM1[1542]<=26'd1970409; ROM2[1542]<=26'd11289329; ROM3[1542]<=26'd9764939; ROM4[1542]<=26'd23472469;
ROM1[1543]<=26'd1963751; ROM2[1543]<=26'd11289061; ROM3[1543]<=26'd9765082; ROM4[1543]<=26'd23472992;
ROM1[1544]<=26'd1948938; ROM2[1544]<=26'd11285433; ROM3[1544]<=26'd9762469; ROM4[1544]<=26'd23468725;
ROM1[1545]<=26'd1943153; ROM2[1545]<=26'd11286259; ROM3[1545]<=26'd9765530; ROM4[1545]<=26'd23468661;
ROM1[1546]<=26'd1942967; ROM2[1546]<=26'd11292400; ROM3[1546]<=26'd9772546; ROM4[1546]<=26'd23472352;
ROM1[1547]<=26'd1944495; ROM2[1547]<=26'd11294088; ROM3[1547]<=26'd9773932; ROM4[1547]<=26'd23472416;
ROM1[1548]<=26'd1947909; ROM2[1548]<=26'd11290200; ROM3[1548]<=26'd9766018; ROM4[1548]<=26'd23469380;
ROM1[1549]<=26'd1967890; ROM2[1549]<=26'd11298070; ROM3[1549]<=26'd9767293; ROM4[1549]<=26'd23476246;
ROM1[1550]<=26'd1989615; ROM2[1550]<=26'd11313512; ROM3[1550]<=26'd9778568; ROM4[1550]<=26'd23489279;
ROM1[1551]<=26'd1978425; ROM2[1551]<=26'd11306126; ROM3[1551]<=26'd9773348; ROM4[1551]<=26'd23482355;
ROM1[1552]<=26'd1957555; ROM2[1552]<=26'd11290687; ROM3[1552]<=26'd9761854; ROM4[1552]<=26'd23466976;
ROM1[1553]<=26'd1949306; ROM2[1553]<=26'd11287125; ROM3[1553]<=26'd9762356; ROM4[1553]<=26'd23464065;
ROM1[1554]<=26'd1939918; ROM2[1554]<=26'd11283692; ROM3[1554]<=26'd9762112; ROM4[1554]<=26'd23462662;
ROM1[1555]<=26'd1934856; ROM2[1555]<=26'd11281006; ROM3[1555]<=26'd9761423; ROM4[1555]<=26'd23460046;
ROM1[1556]<=26'd1942174; ROM2[1556]<=26'd11285188; ROM3[1556]<=26'd9763125; ROM4[1556]<=26'd23462493;
ROM1[1557]<=26'd1946155; ROM2[1557]<=26'd11282017; ROM3[1557]<=26'd9753392; ROM4[1557]<=26'd23457248;
ROM1[1558]<=26'd1951838; ROM2[1558]<=26'd11275923; ROM3[1558]<=26'd9743276; ROM4[1558]<=26'd23450926;
ROM1[1559]<=26'd1957177; ROM2[1559]<=26'd11280928; ROM3[1559]<=26'd9748360; ROM4[1559]<=26'd23456035;
ROM1[1560]<=26'd1960277; ROM2[1560]<=26'd11289720; ROM3[1560]<=26'd9761349; ROM4[1560]<=26'd23467124;
ROM1[1561]<=26'd1959376; ROM2[1561]<=26'd11293683; ROM3[1561]<=26'd9768854; ROM4[1561]<=26'd23473272;
ROM1[1562]<=26'd1949749; ROM2[1562]<=26'd11288803; ROM3[1562]<=26'd9766406; ROM4[1562]<=26'd23469858;
ROM1[1563]<=26'd1940687; ROM2[1563]<=26'd11285265; ROM3[1563]<=26'd9764250; ROM4[1563]<=26'd23465601;
ROM1[1564]<=26'd1933763; ROM2[1564]<=26'd11279400; ROM3[1564]<=26'd9756579; ROM4[1564]<=26'd23457781;
ROM1[1565]<=26'd1937236; ROM2[1565]<=26'd11274606; ROM3[1565]<=26'd9747339; ROM4[1565]<=26'd23452720;
ROM1[1566]<=26'd1958858; ROM2[1566]<=26'd11284845; ROM3[1566]<=26'd9750304; ROM4[1566]<=26'd23459477;
ROM1[1567]<=26'd1971153; ROM2[1567]<=26'd11296032; ROM3[1567]<=26'd9757771; ROM4[1567]<=26'd23468448;
ROM1[1568]<=26'd1961791; ROM2[1568]<=26'd11293020; ROM3[1568]<=26'd9758638; ROM4[1568]<=26'd23467102;
ROM1[1569]<=26'd1951491; ROM2[1569]<=26'd11289780; ROM3[1569]<=26'd9759171; ROM4[1569]<=26'd23464106;
ROM1[1570]<=26'd1952420; ROM2[1570]<=26'd11294003; ROM3[1570]<=26'd9764848; ROM4[1570]<=26'd23467505;
ROM1[1571]<=26'd1944854; ROM2[1571]<=26'd11290574; ROM3[1571]<=26'd9765132; ROM4[1571]<=26'd23465030;
ROM1[1572]<=26'd1938460; ROM2[1572]<=26'd11285724; ROM3[1572]<=26'd9759436; ROM4[1572]<=26'd23459638;
ROM1[1573]<=26'd1949416; ROM2[1573]<=26'd11290146; ROM3[1573]<=26'd9760713; ROM4[1573]<=26'd23463619;
ROM1[1574]<=26'd1956694; ROM2[1574]<=26'd11286573; ROM3[1574]<=26'd9753190; ROM4[1574]<=26'd23459847;
ROM1[1575]<=26'd1950442; ROM2[1575]<=26'd11274378; ROM3[1575]<=26'd9739280; ROM4[1575]<=26'd23448749;
ROM1[1576]<=26'd1952023; ROM2[1576]<=26'd11279240; ROM3[1576]<=26'd9747486; ROM4[1576]<=26'd23454606;
ROM1[1577]<=26'd1952837; ROM2[1577]<=26'd11287245; ROM3[1577]<=26'd9760772; ROM4[1577]<=26'd23463986;
ROM1[1578]<=26'd1950326; ROM2[1578]<=26'd11289915; ROM3[1578]<=26'd9767508; ROM4[1578]<=26'd23469987;
ROM1[1579]<=26'd1949714; ROM2[1579]<=26'd11294392; ROM3[1579]<=26'd9775069; ROM4[1579]<=26'd23475954;
ROM1[1580]<=26'd1947070; ROM2[1580]<=26'd11296213; ROM3[1580]<=26'd9778831; ROM4[1580]<=26'd23475744;
ROM1[1581]<=26'd1951468; ROM2[1581]<=26'd11297063; ROM3[1581]<=26'd9778192; ROM4[1581]<=26'd23476256;
ROM1[1582]<=26'd1962004; ROM2[1582]<=26'd11297382; ROM3[1582]<=26'd9774537; ROM4[1582]<=26'd23476689;
ROM1[1583]<=26'd1965667; ROM2[1583]<=26'd11291404; ROM3[1583]<=26'd9763644; ROM4[1583]<=26'd23470404;
ROM1[1584]<=26'd1963986; ROM2[1584]<=26'd11288656; ROM3[1584]<=26'd9763267; ROM4[1584]<=26'd23471000;
ROM1[1585]<=26'd1956677; ROM2[1585]<=26'd11286829; ROM3[1585]<=26'd9766897; ROM4[1585]<=26'd23469549;
ROM1[1586]<=26'd1950076; ROM2[1586]<=26'd11287933; ROM3[1586]<=26'd9771329; ROM4[1586]<=26'd23470871;
ROM1[1587]<=26'd1960745; ROM2[1587]<=26'd11303870; ROM3[1587]<=26'd9791078; ROM4[1587]<=26'd23487666;
ROM1[1588]<=26'd1959821; ROM2[1588]<=26'd11307141; ROM3[1588]<=26'd9795852; ROM4[1588]<=26'd23490555;
ROM1[1589]<=26'd1949039; ROM2[1589]<=26'd11294886; ROM3[1589]<=26'd9780843; ROM4[1589]<=26'd23477837;
ROM1[1590]<=26'd1951231; ROM2[1590]<=26'd11287944; ROM3[1590]<=26'd9768473; ROM4[1590]<=26'd23468424;
ROM1[1591]<=26'd1964492; ROM2[1591]<=26'd11288247; ROM3[1591]<=26'd9763146; ROM4[1591]<=26'd23469365;
ROM1[1592]<=26'd1971925; ROM2[1592]<=26'd11292316; ROM3[1592]<=26'd9764482; ROM4[1592]<=26'd23472761;
ROM1[1593]<=26'd1965673; ROM2[1593]<=26'd11292136; ROM3[1593]<=26'd9767293; ROM4[1593]<=26'd23473133;
ROM1[1594]<=26'd1958652; ROM2[1594]<=26'd11292810; ROM3[1594]<=26'd9773107; ROM4[1594]<=26'd23473679;
ROM1[1595]<=26'd1953051; ROM2[1595]<=26'd11290379; ROM3[1595]<=26'd9772402; ROM4[1595]<=26'd23471664;
ROM1[1596]<=26'd1944916; ROM2[1596]<=26'd11287458; ROM3[1596]<=26'd9772444; ROM4[1596]<=26'd23471450;
ROM1[1597]<=26'd1944713; ROM2[1597]<=26'd11291071; ROM3[1597]<=26'd9775782; ROM4[1597]<=26'd23472760;
ROM1[1598]<=26'd1951554; ROM2[1598]<=26'd11294183; ROM3[1598]<=26'd9774046; ROM4[1598]<=26'd23473856;
ROM1[1599]<=26'd1962961; ROM2[1599]<=26'd11295883; ROM3[1599]<=26'd9766535; ROM4[1599]<=26'd23470602;
ROM1[1600]<=26'd1969122; ROM2[1600]<=26'd11293823; ROM3[1600]<=26'd9760674; ROM4[1600]<=26'd23466367;
ROM1[1601]<=26'd1964750; ROM2[1601]<=26'd11292119; ROM3[1601]<=26'd9761323; ROM4[1601]<=26'd23465856;
ROM1[1602]<=26'd1960040; ROM2[1602]<=26'd11294312; ROM3[1602]<=26'd9766420; ROM4[1602]<=26'd23468723;
ROM1[1603]<=26'd1961125; ROM2[1603]<=26'd11301252; ROM3[1603]<=26'd9776880; ROM4[1603]<=26'd23476221;
ROM1[1604]<=26'd1954539; ROM2[1604]<=26'd11302024; ROM3[1604]<=26'd9779158; ROM4[1604]<=26'd23477013;
ROM1[1605]<=26'd1938459; ROM2[1605]<=26'd11289141; ROM3[1605]<=26'd9767000; ROM4[1605]<=26'd23463886;
ROM1[1606]<=26'd1936767; ROM2[1606]<=26'd11282348; ROM3[1606]<=26'd9759010; ROM4[1606]<=26'd23455662;
ROM1[1607]<=26'd1945164; ROM2[1607]<=26'd11280951; ROM3[1607]<=26'd9751436; ROM4[1607]<=26'd23453515;
ROM1[1608]<=26'd1960460; ROM2[1608]<=26'd11285758; ROM3[1608]<=26'd9751186; ROM4[1608]<=26'd23457219;
ROM1[1609]<=26'd1976662; ROM2[1609]<=26'd11301757; ROM3[1609]<=26'd9768405; ROM4[1609]<=26'd23473237;
ROM1[1610]<=26'd1967316; ROM2[1610]<=26'd11299119; ROM3[1610]<=26'd9768956; ROM4[1610]<=26'd23472118;
ROM1[1611]<=26'd1948075; ROM2[1611]<=26'd11284385; ROM3[1611]<=26'd9757562; ROM4[1611]<=26'd23456923;
ROM1[1612]<=26'd1939878; ROM2[1612]<=26'd11279498; ROM3[1612]<=26'd9754567; ROM4[1612]<=26'd23452570;
ROM1[1613]<=26'd1932086; ROM2[1613]<=26'd11276144; ROM3[1613]<=26'd9752155; ROM4[1613]<=26'd23450792;
ROM1[1614]<=26'd1934643; ROM2[1614]<=26'd11277583; ROM3[1614]<=26'd9750745; ROM4[1614]<=26'd23451104;
ROM1[1615]<=26'd1944219; ROM2[1615]<=26'd11281563; ROM3[1615]<=26'd9751881; ROM4[1615]<=26'd23452661;
ROM1[1616]<=26'd1954565; ROM2[1616]<=26'd11283560; ROM3[1616]<=26'd9747001; ROM4[1616]<=26'd23452256;
ROM1[1617]<=26'd1959174; ROM2[1617]<=26'd11285613; ROM3[1617]<=26'd9744857; ROM4[1617]<=26'd23453048;
ROM1[1618]<=26'd1950900; ROM2[1618]<=26'd11281311; ROM3[1618]<=26'd9742884; ROM4[1618]<=26'd23450875;
ROM1[1619]<=26'd1951834; ROM2[1619]<=26'd11288257; ROM3[1619]<=26'd9754259; ROM4[1619]<=26'd23458877;
ROM1[1620]<=26'd1951146; ROM2[1620]<=26'd11291108; ROM3[1620]<=26'd9761669; ROM4[1620]<=26'd23462348;
ROM1[1621]<=26'd1935343; ROM2[1621]<=26'd11279702; ROM3[1621]<=26'd9755401; ROM4[1621]<=26'd23451151;
ROM1[1622]<=26'd1929862; ROM2[1622]<=26'd11274992; ROM3[1622]<=26'd9754952; ROM4[1622]<=26'd23446766;
ROM1[1623]<=26'd1930778; ROM2[1623]<=26'd11269996; ROM3[1623]<=26'd9747644; ROM4[1623]<=26'd23442496;
ROM1[1624]<=26'd1941588; ROM2[1624]<=26'd11269128; ROM3[1624]<=26'd9741251; ROM4[1624]<=26'd23439548;
ROM1[1625]<=26'd1953143; ROM2[1625]<=26'd11272910; ROM3[1625]<=26'd9741537; ROM4[1625]<=26'd23443933;
ROM1[1626]<=26'd1950212; ROM2[1626]<=26'd11275117; ROM3[1626]<=26'd9746697; ROM4[1626]<=26'd23447373;
ROM1[1627]<=26'd1942440; ROM2[1627]<=26'd11276822; ROM3[1627]<=26'd9750512; ROM4[1627]<=26'd23448347;
ROM1[1628]<=26'd1939432; ROM2[1628]<=26'd11280192; ROM3[1628]<=26'd9756003; ROM4[1628]<=26'd23453253;
ROM1[1629]<=26'd1934627; ROM2[1629]<=26'd11281362; ROM3[1629]<=26'd9761595; ROM4[1629]<=26'd23455266;
ROM1[1630]<=26'd1934911; ROM2[1630]<=26'd11285112; ROM3[1630]<=26'd9763860; ROM4[1630]<=26'd23457741;
ROM1[1631]<=26'd1946451; ROM2[1631]<=26'd11293023; ROM3[1631]<=26'd9768234; ROM4[1631]<=26'd23463854;
ROM1[1632]<=26'd1956841; ROM2[1632]<=26'd11292244; ROM3[1632]<=26'd9763003; ROM4[1632]<=26'd23463363;
ROM1[1633]<=26'd1965430; ROM2[1633]<=26'd11291354; ROM3[1633]<=26'd9757259; ROM4[1633]<=26'd23463653;
ROM1[1634]<=26'd1964537; ROM2[1634]<=26'd11291324; ROM3[1634]<=26'd9758103; ROM4[1634]<=26'd23463469;
ROM1[1635]<=26'd1958238; ROM2[1635]<=26'd11289193; ROM3[1635]<=26'd9760716; ROM4[1635]<=26'd23463141;
ROM1[1636]<=26'd1956822; ROM2[1636]<=26'd11295736; ROM3[1636]<=26'd9769823; ROM4[1636]<=26'd23470429;
ROM1[1637]<=26'd1958472; ROM2[1637]<=26'd11303939; ROM3[1637]<=26'd9778113; ROM4[1637]<=26'd23477429;
ROM1[1638]<=26'd1953150; ROM2[1638]<=26'd11301973; ROM3[1638]<=26'd9778948; ROM4[1638]<=26'd23476677;
ROM1[1639]<=26'd1950028; ROM2[1639]<=26'd11296876; ROM3[1639]<=26'd9774132; ROM4[1639]<=26'd23471822;
ROM1[1640]<=26'd1956704; ROM2[1640]<=26'd11293881; ROM3[1640]<=26'd9767201; ROM4[1640]<=26'd23466566;
ROM1[1641]<=26'd1971286; ROM2[1641]<=26'd11297415; ROM3[1641]<=26'd9763312; ROM4[1641]<=26'd23467237;
ROM1[1642]<=26'd1982196; ROM2[1642]<=26'd11305287; ROM3[1642]<=26'd9767207; ROM4[1642]<=26'd23474767;
ROM1[1643]<=26'd1976363; ROM2[1643]<=26'd11303333; ROM3[1643]<=26'd9769175; ROM4[1643]<=26'd23475084;
ROM1[1644]<=26'd1964330; ROM2[1644]<=26'd11297953; ROM3[1644]<=26'd9770885; ROM4[1644]<=26'd23471999;
ROM1[1645]<=26'd1955113; ROM2[1645]<=26'd11293487; ROM3[1645]<=26'd9772601; ROM4[1645]<=26'd23470907;
ROM1[1646]<=26'd1948052; ROM2[1646]<=26'd11291899; ROM3[1646]<=26'd9772647; ROM4[1646]<=26'd23469605;
ROM1[1647]<=26'd1952284; ROM2[1647]<=26'd11294253; ROM3[1647]<=26'd9774684; ROM4[1647]<=26'd23471560;
ROM1[1648]<=26'd1961215; ROM2[1648]<=26'd11294942; ROM3[1648]<=26'd9771824; ROM4[1648]<=26'd23471757;
ROM1[1649]<=26'd1979766; ROM2[1649]<=26'd11300632; ROM3[1649]<=26'd9768996; ROM4[1649]<=26'd23476571;
ROM1[1650]<=26'd1995138; ROM2[1650]<=26'd11307257; ROM3[1650]<=26'd9773167; ROM4[1650]<=26'd23484235;
ROM1[1651]<=26'd1990428; ROM2[1651]<=26'd11308307; ROM3[1651]<=26'd9776059; ROM4[1651]<=26'd23485923;
ROM1[1652]<=26'd1977801; ROM2[1652]<=26'd11301977; ROM3[1652]<=26'd9773920; ROM4[1652]<=26'd23482837;
ROM1[1653]<=26'd1970708; ROM2[1653]<=26'd11298716; ROM3[1653]<=26'd9775411; ROM4[1653]<=26'd23482059;
ROM1[1654]<=26'd1957005; ROM2[1654]<=26'd11290939; ROM3[1654]<=26'd9770815; ROM4[1654]<=26'd23475123;
ROM1[1655]<=26'd1945391; ROM2[1655]<=26'd11282395; ROM3[1655]<=26'd9762802; ROM4[1655]<=26'd23465630;
ROM1[1656]<=26'd1954748; ROM2[1656]<=26'd11289466; ROM3[1656]<=26'd9765331; ROM4[1656]<=26'd23468539;
ROM1[1657]<=26'd1967446; ROM2[1657]<=26'd11292257; ROM3[1657]<=26'd9762056; ROM4[1657]<=26'd23467939;
ROM1[1658]<=26'd1974978; ROM2[1658]<=26'd11289664; ROM3[1658]<=26'd9754105; ROM4[1658]<=26'd23464053;
ROM1[1659]<=26'd1974906; ROM2[1659]<=26'd11291165; ROM3[1659]<=26'd9755679; ROM4[1659]<=26'd23466469;
ROM1[1660]<=26'd1970542; ROM2[1660]<=26'd11293564; ROM3[1660]<=26'd9760790; ROM4[1660]<=26'd23469763;
ROM1[1661]<=26'd1963406; ROM2[1661]<=26'd11291278; ROM3[1661]<=26'd9764388; ROM4[1661]<=26'd23469056;
ROM1[1662]<=26'd1953507; ROM2[1662]<=26'd11287241; ROM3[1662]<=26'd9762861; ROM4[1662]<=26'd23466158;
ROM1[1663]<=26'd1945910; ROM2[1663]<=26'd11287158; ROM3[1663]<=26'd9764867; ROM4[1663]<=26'd23466123;
ROM1[1664]<=26'd1947113; ROM2[1664]<=26'd11289222; ROM3[1664]<=26'd9766763; ROM4[1664]<=26'd23469353;
ROM1[1665]<=26'd1956310; ROM2[1665]<=26'd11291508; ROM3[1665]<=26'd9763977; ROM4[1665]<=26'd23470429;
ROM1[1666]<=26'd1969963; ROM2[1666]<=26'd11292711; ROM3[1666]<=26'd9759494; ROM4[1666]<=26'd23470194;
ROM1[1667]<=26'd1973422; ROM2[1667]<=26'd11291735; ROM3[1667]<=26'd9756697; ROM4[1667]<=26'd23470439;
ROM1[1668]<=26'd1961026; ROM2[1668]<=26'd11282993; ROM3[1668]<=26'd9752944; ROM4[1668]<=26'd23463808;
ROM1[1669]<=26'd1950126; ROM2[1669]<=26'd11278677; ROM3[1669]<=26'd9751510; ROM4[1669]<=26'd23460187;
ROM1[1670]<=26'd1946625; ROM2[1670]<=26'd11282484; ROM3[1670]<=26'd9757058; ROM4[1670]<=26'd23463357;
ROM1[1671]<=26'd1940312; ROM2[1671]<=26'd11282023; ROM3[1671]<=26'd9760294; ROM4[1671]<=26'd23462791;
ROM1[1672]<=26'd1937404; ROM2[1672]<=26'd11281004; ROM3[1672]<=26'd9757728; ROM4[1672]<=26'd23459333;
ROM1[1673]<=26'd1946809; ROM2[1673]<=26'd11285209; ROM3[1673]<=26'd9757329; ROM4[1673]<=26'd23460472;
ROM1[1674]<=26'd1960905; ROM2[1674]<=26'd11287133; ROM3[1674]<=26'd9753136; ROM4[1674]<=26'd23460676;
ROM1[1675]<=26'd1964793; ROM2[1675]<=26'd11284791; ROM3[1675]<=26'd9746826; ROM4[1675]<=26'd23458109;
ROM1[1676]<=26'd1956169; ROM2[1676]<=26'd11279099; ROM3[1676]<=26'd9743533; ROM4[1676]<=26'd23453273;
ROM1[1677]<=26'd1944733; ROM2[1677]<=26'd11274491; ROM3[1677]<=26'd9742389; ROM4[1677]<=26'd23448589;
ROM1[1678]<=26'd1936962; ROM2[1678]<=26'd11272484; ROM3[1678]<=26'd9742719; ROM4[1678]<=26'd23446123;
ROM1[1679]<=26'd1934216; ROM2[1679]<=26'd11273549; ROM3[1679]<=26'd9746918; ROM4[1679]<=26'd23447157;
ROM1[1680]<=26'd1935039; ROM2[1680]<=26'd11278465; ROM3[1680]<=26'd9750403; ROM4[1680]<=26'd23451559;
ROM1[1681]<=26'd1938403; ROM2[1681]<=26'd11279598; ROM3[1681]<=26'd9748333; ROM4[1681]<=26'd23452771;
ROM1[1682]<=26'd1948472; ROM2[1682]<=26'd11278572; ROM3[1682]<=26'd9742715; ROM4[1682]<=26'd23450741;
ROM1[1683]<=26'd1956553; ROM2[1683]<=26'd11277215; ROM3[1683]<=26'd9735004; ROM4[1683]<=26'd23448376;
ROM1[1684]<=26'd1955639; ROM2[1684]<=26'd11277386; ROM3[1684]<=26'd9735578; ROM4[1684]<=26'd23447608;
ROM1[1685]<=26'd1948515; ROM2[1685]<=26'd11275122; ROM3[1685]<=26'd9738564; ROM4[1685]<=26'd23446150;
ROM1[1686]<=26'd1940738; ROM2[1686]<=26'd11273832; ROM3[1686]<=26'd9742266; ROM4[1686]<=26'd23446785;
ROM1[1687]<=26'd1934837; ROM2[1687]<=26'd11274791; ROM3[1687]<=26'd9743911; ROM4[1687]<=26'd23447747;
ROM1[1688]<=26'd1934418; ROM2[1688]<=26'd11277397; ROM3[1688]<=26'd9747490; ROM4[1688]<=26'd23450436;
ROM1[1689]<=26'd1946051; ROM2[1689]<=26'd11285887; ROM3[1689]<=26'd9754589; ROM4[1689]<=26'd23457624;
ROM1[1690]<=26'd1959109; ROM2[1690]<=26'd11290962; ROM3[1690]<=26'd9755545; ROM4[1690]<=26'd23461650;
ROM1[1691]<=26'd1968099; ROM2[1691]<=26'd11289733; ROM3[1691]<=26'd9748941; ROM4[1691]<=26'd23459715;
ROM1[1692]<=26'd1964616; ROM2[1692]<=26'd11285123; ROM3[1692]<=26'd9743055; ROM4[1692]<=26'd23454595;
ROM1[1693]<=26'd1953600; ROM2[1693]<=26'd11279534; ROM3[1693]<=26'd9741068; ROM4[1693]<=26'd23450246;
ROM1[1694]<=26'd1942934; ROM2[1694]<=26'd11273791; ROM3[1694]<=26'd9740743; ROM4[1694]<=26'd23447070;
ROM1[1695]<=26'd1939471; ROM2[1695]<=26'd11272461; ROM3[1695]<=26'd9743915; ROM4[1695]<=26'd23447530;
ROM1[1696]<=26'd1938590; ROM2[1696]<=26'd11276527; ROM3[1696]<=26'd9752371; ROM4[1696]<=26'd23453961;
ROM1[1697]<=26'd1944252; ROM2[1697]<=26'd11283629; ROM3[1697]<=26'd9759823; ROM4[1697]<=26'd23461741;
ROM1[1698]<=26'd1953108; ROM2[1698]<=26'd11286820; ROM3[1698]<=26'd9759168; ROM4[1698]<=26'd23463444;
ROM1[1699]<=26'd1966779; ROM2[1699]<=26'd11290622; ROM3[1699]<=26'd9755664; ROM4[1699]<=26'd23464901;
ROM1[1700]<=26'd1969036; ROM2[1700]<=26'd11286666; ROM3[1700]<=26'd9748455; ROM4[1700]<=26'd23460453;
ROM1[1701]<=26'd1952179; ROM2[1701]<=26'd11273085; ROM3[1701]<=26'd9739570; ROM4[1701]<=26'd23448991;
ROM1[1702]<=26'd1946117; ROM2[1702]<=26'd11274437; ROM3[1702]<=26'd9743008; ROM4[1702]<=26'd23450402;
ROM1[1703]<=26'd1948653; ROM2[1703]<=26'd11281696; ROM3[1703]<=26'd9753734; ROM4[1703]<=26'd23457675;
ROM1[1704]<=26'd1948272; ROM2[1704]<=26'd11285197; ROM3[1704]<=26'd9761462; ROM4[1704]<=26'd23462893;
ROM1[1705]<=26'd1945730; ROM2[1705]<=26'd11285860; ROM3[1705]<=26'd9763811; ROM4[1705]<=26'd23463817;
ROM1[1706]<=26'd1947342; ROM2[1706]<=26'd11285275; ROM3[1706]<=26'd9763996; ROM4[1706]<=26'd23463195;
ROM1[1707]<=26'd1960710; ROM2[1707]<=26'd11287233; ROM3[1707]<=26'd9760323; ROM4[1707]<=26'd23464713;
ROM1[1708]<=26'd1971222; ROM2[1708]<=26'd11287517; ROM3[1708]<=26'd9753442; ROM4[1708]<=26'd23463851;
ROM1[1709]<=26'd1969047; ROM2[1709]<=26'd11287992; ROM3[1709]<=26'd9753866; ROM4[1709]<=26'd23464451;
ROM1[1710]<=26'd1963577; ROM2[1710]<=26'd11289342; ROM3[1710]<=26'd9758643; ROM4[1710]<=26'd23467157;
ROM1[1711]<=26'd1959097; ROM2[1711]<=26'd11290736; ROM3[1711]<=26'd9764126; ROM4[1711]<=26'd23469459;
ROM1[1712]<=26'd1955903; ROM2[1712]<=26'd11294953; ROM3[1712]<=26'd9771038; ROM4[1712]<=26'd23473014;
ROM1[1713]<=26'd1945987; ROM2[1713]<=26'd11289551; ROM3[1713]<=26'd9767687; ROM4[1713]<=26'd23466363;
ROM1[1714]<=26'd1947200; ROM2[1714]<=26'd11287042; ROM3[1714]<=26'd9763885; ROM4[1714]<=26'd23463800;
ROM1[1715]<=26'd1957854; ROM2[1715]<=26'd11289672; ROM3[1715]<=26'd9762066; ROM4[1715]<=26'd23464960;
ROM1[1716]<=26'd1971600; ROM2[1716]<=26'd11290791; ROM3[1716]<=26'd9758373; ROM4[1716]<=26'd23464867;
ROM1[1717]<=26'd1976192; ROM2[1717]<=26'd11293760; ROM3[1717]<=26'd9757703; ROM4[1717]<=26'd23467401;
ROM1[1718]<=26'd1965981; ROM2[1718]<=26'd11290534; ROM3[1718]<=26'd9758799; ROM4[1718]<=26'd23465900;
ROM1[1719]<=26'd1957364; ROM2[1719]<=26'd11287707; ROM3[1719]<=26'd9761047; ROM4[1719]<=26'd23465509;
ROM1[1720]<=26'd1954915; ROM2[1720]<=26'd11287758; ROM3[1720]<=26'd9763639; ROM4[1720]<=26'd23467058;
ROM1[1721]<=26'd1951653; ROM2[1721]<=26'd11287077; ROM3[1721]<=26'd9768904; ROM4[1721]<=26'd23470132;
ROM1[1722]<=26'd1954516; ROM2[1722]<=26'd11290850; ROM3[1722]<=26'd9771398; ROM4[1722]<=26'd23472680;
ROM1[1723]<=26'd1961866; ROM2[1723]<=26'd11293470; ROM3[1723]<=26'd9769997; ROM4[1723]<=26'd23473662;
ROM1[1724]<=26'd1972759; ROM2[1724]<=26'd11293970; ROM3[1724]<=26'd9765111; ROM4[1724]<=26'd23471768;
ROM1[1725]<=26'd1980683; ROM2[1725]<=26'd11295563; ROM3[1725]<=26'd9763991; ROM4[1725]<=26'd23472919;
ROM1[1726]<=26'd1978055; ROM2[1726]<=26'd11296698; ROM3[1726]<=26'd9767343; ROM4[1726]<=26'd23474912;
ROM1[1727]<=26'd1967296; ROM2[1727]<=26'd11293364; ROM3[1727]<=26'd9767282; ROM4[1727]<=26'd23471493;
ROM1[1728]<=26'd1961638; ROM2[1728]<=26'd11292573; ROM3[1728]<=26'd9771197; ROM4[1728]<=26'd23473435;
ROM1[1729]<=26'd1956845; ROM2[1729]<=26'd11293134; ROM3[1729]<=26'd9772796; ROM4[1729]<=26'd23472497;
ROM1[1730]<=26'd1950049; ROM2[1730]<=26'd11288554; ROM3[1730]<=26'd9767350; ROM4[1730]<=26'd23466939;
ROM1[1731]<=26'd1954546; ROM2[1731]<=26'd11288585; ROM3[1731]<=26'd9767854; ROM4[1731]<=26'd23469229;
ROM1[1732]<=26'd1965701; ROM2[1732]<=26'd11289765; ROM3[1732]<=26'd9763167; ROM4[1732]<=26'd23469041;
ROM1[1733]<=26'd1978637; ROM2[1733]<=26'd11294500; ROM3[1733]<=26'd9759502; ROM4[1733]<=26'd23472099;
ROM1[1734]<=26'd1978886; ROM2[1734]<=26'd11295691; ROM3[1734]<=26'd9759901; ROM4[1734]<=26'd23472089;
ROM1[1735]<=26'd1969866; ROM2[1735]<=26'd11292052; ROM3[1735]<=26'd9759326; ROM4[1735]<=26'd23468264;
ROM1[1736]<=26'd1963030; ROM2[1736]<=26'd11290971; ROM3[1736]<=26'd9763144; ROM4[1736]<=26'd23468395;
ROM1[1737]<=26'd1961388; ROM2[1737]<=26'd11294110; ROM3[1737]<=26'd9767286; ROM4[1737]<=26'd23470998;
ROM1[1738]<=26'd1957666; ROM2[1738]<=26'd11294068; ROM3[1738]<=26'd9769454; ROM4[1738]<=26'd23472722;
ROM1[1739]<=26'd1954623; ROM2[1739]<=26'd11291021; ROM3[1739]<=26'd9765421; ROM4[1739]<=26'd23468040;
ROM1[1740]<=26'd1965056; ROM2[1740]<=26'd11294216; ROM3[1740]<=26'd9761485; ROM4[1740]<=26'd23468107;
ROM1[1741]<=26'd1976214; ROM2[1741]<=26'd11294450; ROM3[1741]<=26'd9755576; ROM4[1741]<=26'd23466637;
ROM1[1742]<=26'd1974562; ROM2[1742]<=26'd11291139; ROM3[1742]<=26'd9749846; ROM4[1742]<=26'd23461470;
ROM1[1743]<=26'd1968230; ROM2[1743]<=26'd11290735; ROM3[1743]<=26'd9751989; ROM4[1743]<=26'd23462472;
ROM1[1744]<=26'd1959645; ROM2[1744]<=26'd11290983; ROM3[1744]<=26'd9755869; ROM4[1744]<=26'd23462563;
ROM1[1745]<=26'd1956641; ROM2[1745]<=26'd11292508; ROM3[1745]<=26'd9761088; ROM4[1745]<=26'd23465304;
ROM1[1746]<=26'd1960914; ROM2[1746]<=26'd11303100; ROM3[1746]<=26'd9775591; ROM4[1746]<=26'd23479112;
ROM1[1747]<=26'd1970257; ROM2[1747]<=26'd11313724; ROM3[1747]<=26'd9785070; ROM4[1747]<=26'd23487466;
ROM1[1748]<=26'd1966906; ROM2[1748]<=26'd11305049; ROM3[1748]<=26'd9770137; ROM4[1748]<=26'd23475180;
ROM1[1749]<=26'd1960582; ROM2[1749]<=26'd11288628; ROM3[1749]<=26'd9747335; ROM4[1749]<=26'd23457624;
ROM1[1750]<=26'd1958814; ROM2[1750]<=26'd11280612; ROM3[1750]<=26'd9738711; ROM4[1750]<=26'd23450671;
ROM1[1751]<=26'd1952428; ROM2[1751]<=26'd11276210; ROM3[1751]<=26'd9739556; ROM4[1751]<=26'd23449271;
ROM1[1752]<=26'd1950856; ROM2[1752]<=26'd11280735; ROM3[1752]<=26'd9750679; ROM4[1752]<=26'd23455267;
ROM1[1753]<=26'd1948601; ROM2[1753]<=26'd11284469; ROM3[1753]<=26'd9758988; ROM4[1753]<=26'd23460438;
ROM1[1754]<=26'd1938684; ROM2[1754]<=26'd11280025; ROM3[1754]<=26'd9757816; ROM4[1754]<=26'd23455941;
ROM1[1755]<=26'd1928722; ROM2[1755]<=26'd11275078; ROM3[1755]<=26'd9753344; ROM4[1755]<=26'd23450286;
ROM1[1756]<=26'd1930635; ROM2[1756]<=26'd11274277; ROM3[1756]<=26'd9751587; ROM4[1756]<=26'd23450672;
ROM1[1757]<=26'd1944610; ROM2[1757]<=26'd11278759; ROM3[1757]<=26'd9752723; ROM4[1757]<=26'd23454074;
ROM1[1758]<=26'd1953679; ROM2[1758]<=26'd11278708; ROM3[1758]<=26'd9746738; ROM4[1758]<=26'd23451925;
ROM1[1759]<=26'd1951818; ROM2[1759]<=26'd11277265; ROM3[1759]<=26'd9742746; ROM4[1759]<=26'd23450228;
ROM1[1760]<=26'd1954884; ROM2[1760]<=26'd11282483; ROM3[1760]<=26'd9753280; ROM4[1760]<=26'd23457962;
ROM1[1761]<=26'd1953194; ROM2[1761]<=26'd11284809; ROM3[1761]<=26'd9760236; ROM4[1761]<=26'd23461166;
ROM1[1762]<=26'd1947089; ROM2[1762]<=26'd11283467; ROM3[1762]<=26'd9760104; ROM4[1762]<=26'd23459412;
ROM1[1763]<=26'd1944007; ROM2[1763]<=26'd11285321; ROM3[1763]<=26'd9763285; ROM4[1763]<=26'd23460728;
ROM1[1764]<=26'd1945527; ROM2[1764]<=26'd11287713; ROM3[1764]<=26'd9762089; ROM4[1764]<=26'd23461592;
ROM1[1765]<=26'd1955977; ROM2[1765]<=26'd11288643; ROM3[1765]<=26'd9756652; ROM4[1765]<=26'd23460888;
ROM1[1766]<=26'd1969416; ROM2[1766]<=26'd11290060; ROM3[1766]<=26'd9752775; ROM4[1766]<=26'd23461482;
ROM1[1767]<=26'd1969779; ROM2[1767]<=26'd11287997; ROM3[1767]<=26'd9750997; ROM4[1767]<=26'd23459484;
ROM1[1768]<=26'd1956208; ROM2[1768]<=26'd11279441; ROM3[1768]<=26'd9746436; ROM4[1768]<=26'd23452593;
ROM1[1769]<=26'd1948270; ROM2[1769]<=26'd11277012; ROM3[1769]<=26'd9748503; ROM4[1769]<=26'd23451680;
ROM1[1770]<=26'd1947328; ROM2[1770]<=26'd11280455; ROM3[1770]<=26'd9754744; ROM4[1770]<=26'd23455234;
ROM1[1771]<=26'd1947197; ROM2[1771]<=26'd11284125; ROM3[1771]<=26'd9760766; ROM4[1771]<=26'd23461062;
ROM1[1772]<=26'd1949940; ROM2[1772]<=26'd11287617; ROM3[1772]<=26'd9762098; ROM4[1772]<=26'd23464758;
ROM1[1773]<=26'd1959407; ROM2[1773]<=26'd11291689; ROM3[1773]<=26'd9762873; ROM4[1773]<=26'd23467151;
ROM1[1774]<=26'd1973112; ROM2[1774]<=26'd11293671; ROM3[1774]<=26'd9758947; ROM4[1774]<=26'd23467765;
ROM1[1775]<=26'd1978360; ROM2[1775]<=26'd11293920; ROM3[1775]<=26'd9754445; ROM4[1775]<=26'd23466825;
ROM1[1776]<=26'd1976251; ROM2[1776]<=26'd11296870; ROM3[1776]<=26'd9757798; ROM4[1776]<=26'd23468611;
ROM1[1777]<=26'd1968972; ROM2[1777]<=26'd11297636; ROM3[1777]<=26'd9759701; ROM4[1777]<=26'd23470152;
ROM1[1778]<=26'd1964200; ROM2[1778]<=26'd11298991; ROM3[1778]<=26'd9762972; ROM4[1778]<=26'd23472355;
ROM1[1779]<=26'd1958435; ROM2[1779]<=26'd11299059; ROM3[1779]<=26'd9768009; ROM4[1779]<=26'd23474075;
ROM1[1780]<=26'd1951911; ROM2[1780]<=26'd11295534; ROM3[1780]<=26'd9766768; ROM4[1780]<=26'd23470854;
ROM1[1781]<=26'd1957438; ROM2[1781]<=26'd11296589; ROM3[1781]<=26'd9767483; ROM4[1781]<=26'd23471985;
ROM1[1782]<=26'd1973506; ROM2[1782]<=26'd11301937; ROM3[1782]<=26'd9766692; ROM4[1782]<=26'd23475496;
ROM1[1783]<=26'd1980887; ROM2[1783]<=26'd11298143; ROM3[1783]<=26'd9757005; ROM4[1783]<=26'd23470851;
ROM1[1784]<=26'd1976171; ROM2[1784]<=26'd11294020; ROM3[1784]<=26'd9754217; ROM4[1784]<=26'd23467605;
ROM1[1785]<=26'd1969741; ROM2[1785]<=26'd11295575; ROM3[1785]<=26'd9759461; ROM4[1785]<=26'd23470888;
ROM1[1786]<=26'd1963618; ROM2[1786]<=26'd11294695; ROM3[1786]<=26'd9764992; ROM4[1786]<=26'd23472697;
ROM1[1787]<=26'd1963148; ROM2[1787]<=26'd11299407; ROM3[1787]<=26'd9772898; ROM4[1787]<=26'd23476434;
ROM1[1788]<=26'd1957136; ROM2[1788]<=26'd11297428; ROM3[1788]<=26'd9772705; ROM4[1788]<=26'd23474646;
ROM1[1789]<=26'd1951248; ROM2[1789]<=26'd11290373; ROM3[1789]<=26'd9766292; ROM4[1789]<=26'd23466587;
ROM1[1790]<=26'd1964057; ROM2[1790]<=26'd11294899; ROM3[1790]<=26'd9766069; ROM4[1790]<=26'd23468450;
ROM1[1791]<=26'd1981169; ROM2[1791]<=26'd11301052; ROM3[1791]<=26'd9762804; ROM4[1791]<=26'd23473280;
ROM1[1792]<=26'd1973705; ROM2[1792]<=26'd11294499; ROM3[1792]<=26'd9752560; ROM4[1792]<=26'd23464938;
ROM1[1793]<=26'd1960825; ROM2[1793]<=26'd11286911; ROM3[1793]<=26'd9747362; ROM4[1793]<=26'd23456481;
ROM1[1794]<=26'd1951539; ROM2[1794]<=26'd11283283; ROM3[1794]<=26'd9747954; ROM4[1794]<=26'd23453856;
ROM1[1795]<=26'd1943142; ROM2[1795]<=26'd11279800; ROM3[1795]<=26'd9747572; ROM4[1795]<=26'd23450246;
ROM1[1796]<=26'd1943710; ROM2[1796]<=26'd11284960; ROM3[1796]<=26'd9754439; ROM4[1796]<=26'd23457359;
ROM1[1797]<=26'd1945179; ROM2[1797]<=26'd11287597; ROM3[1797]<=26'd9753437; ROM4[1797]<=26'd23459378;
ROM1[1798]<=26'd1946098; ROM2[1798]<=26'd11283423; ROM3[1798]<=26'd9743194; ROM4[1798]<=26'd23453817;
ROM1[1799]<=26'd1958889; ROM2[1799]<=26'd11284128; ROM3[1799]<=26'd9739188; ROM4[1799]<=26'd23454080;
ROM1[1800]<=26'd1968991; ROM2[1800]<=26'd11285962; ROM3[1800]<=26'd9739001; ROM4[1800]<=26'd23455195;
ROM1[1801]<=26'd1968199; ROM2[1801]<=26'd11286121; ROM3[1801]<=26'd9742235; ROM4[1801]<=26'd23457120;
ROM1[1802]<=26'd1958887; ROM2[1802]<=26'd11282674; ROM3[1802]<=26'd9743437; ROM4[1802]<=26'd23455960;
ROM1[1803]<=26'd1951932; ROM2[1803]<=26'd11281204; ROM3[1803]<=26'd9745842; ROM4[1803]<=26'd23455727;
ROM1[1804]<=26'd1948346; ROM2[1804]<=26'd11284874; ROM3[1804]<=26'd9751939; ROM4[1804]<=26'd23460298;
ROM1[1805]<=26'd1946439; ROM2[1805]<=26'd11288249; ROM3[1805]<=26'd9755389; ROM4[1805]<=26'd23463960;
ROM1[1806]<=26'd1958327; ROM2[1806]<=26'd11297554; ROM3[1806]<=26'd9760437; ROM4[1806]<=26'd23470614;
ROM1[1807]<=26'd1972629; ROM2[1807]<=26'd11301349; ROM3[1807]<=26'd9757746; ROM4[1807]<=26'd23472320;
ROM1[1808]<=26'd1972465; ROM2[1808]<=26'd11290256; ROM3[1808]<=26'd9742867; ROM4[1808]<=26'd23461559;
ROM1[1809]<=26'd1964642; ROM2[1809]<=26'd11285035; ROM3[1809]<=26'd9738719; ROM4[1809]<=26'd23455616;
ROM1[1810]<=26'd1955918; ROM2[1810]<=26'd11283713; ROM3[1810]<=26'd9740800; ROM4[1810]<=26'd23454488;
ROM1[1811]<=26'd1946775; ROM2[1811]<=26'd11280867; ROM3[1811]<=26'd9739850; ROM4[1811]<=26'd23451005;
ROM1[1812]<=26'd1944388; ROM2[1812]<=26'd11283921; ROM3[1812]<=26'd9746018; ROM4[1812]<=26'd23454166;
ROM1[1813]<=26'd1942160; ROM2[1813]<=26'd11285078; ROM3[1813]<=26'd9751405; ROM4[1813]<=26'd23456509;
ROM1[1814]<=26'd1944581; ROM2[1814]<=26'd11286098; ROM3[1814]<=26'd9750895; ROM4[1814]<=26'd23457453;
ROM1[1815]<=26'd1960300; ROM2[1815]<=26'd11296232; ROM3[1815]<=26'd9753693; ROM4[1815]<=26'd23464544;
ROM1[1816]<=26'd1980214; ROM2[1816]<=26'd11304447; ROM3[1816]<=26'd9753651; ROM4[1816]<=26'd23470599;
ROM1[1817]<=26'd1981480; ROM2[1817]<=26'd11302621; ROM3[1817]<=26'd9751932; ROM4[1817]<=26'd23470016;
ROM1[1818]<=26'd1963720; ROM2[1818]<=26'd11291938; ROM3[1818]<=26'd9747390; ROM4[1818]<=26'd23461821;
ROM1[1819]<=26'd1947860; ROM2[1819]<=26'd11282008; ROM3[1819]<=26'd9746467; ROM4[1819]<=26'd23455749;
ROM1[1820]<=26'd1943599; ROM2[1820]<=26'd11282487; ROM3[1820]<=26'd9750479; ROM4[1820]<=26'd23457405;
ROM1[1821]<=26'd1938597; ROM2[1821]<=26'd11283012; ROM3[1821]<=26'd9754167; ROM4[1821]<=26'd23458351;
ROM1[1822]<=26'd1942388; ROM2[1822]<=26'd11286091; ROM3[1822]<=26'd9758831; ROM4[1822]<=26'd23461831;
ROM1[1823]<=26'd1949832; ROM2[1823]<=26'd11286775; ROM3[1823]<=26'd9756635; ROM4[1823]<=26'd23463256;
ROM1[1824]<=26'd1961193; ROM2[1824]<=26'd11286203; ROM3[1824]<=26'd9750483; ROM4[1824]<=26'd23461779;
ROM1[1825]<=26'd1971037; ROM2[1825]<=26'd11290972; ROM3[1825]<=26'd9749325; ROM4[1825]<=26'd23465519;
ROM1[1826]<=26'd1967332; ROM2[1826]<=26'd11291765; ROM3[1826]<=26'd9750821; ROM4[1826]<=26'd23466365;
ROM1[1827]<=26'd1957893; ROM2[1827]<=26'd11288633; ROM3[1827]<=26'd9753318; ROM4[1827]<=26'd23463859;
ROM1[1828]<=26'd1954489; ROM2[1828]<=26'd11291938; ROM3[1828]<=26'd9759670; ROM4[1828]<=26'd23466299;
ROM1[1829]<=26'd1951856; ROM2[1829]<=26'd11295799; ROM3[1829]<=26'd9764993; ROM4[1829]<=26'd23468890;
ROM1[1830]<=26'd1943403; ROM2[1830]<=26'd11290713; ROM3[1830]<=26'd9763388; ROM4[1830]<=26'd23464909;
ROM1[1831]<=26'd1945549; ROM2[1831]<=26'd11288347; ROM3[1831]<=26'd9759728; ROM4[1831]<=26'd23463132;
ROM1[1832]<=26'd1956154; ROM2[1832]<=26'd11288606; ROM3[1832]<=26'd9755500; ROM4[1832]<=26'd23461470;
ROM1[1833]<=26'd1962464; ROM2[1833]<=26'd11285160; ROM3[1833]<=26'd9749319; ROM4[1833]<=26'd23458742;
ROM1[1834]<=26'd1964077; ROM2[1834]<=26'd11285384; ROM3[1834]<=26'd9749113; ROM4[1834]<=26'd23460960;
ROM1[1835]<=26'd1960879; ROM2[1835]<=26'd11287110; ROM3[1835]<=26'd9753126; ROM4[1835]<=26'd23463123;
ROM1[1836]<=26'd1954592; ROM2[1836]<=26'd11286479; ROM3[1836]<=26'd9758328; ROM4[1836]<=26'd23464075;
ROM1[1837]<=26'd1948415; ROM2[1837]<=26'd11286441; ROM3[1837]<=26'd9761781; ROM4[1837]<=26'd23465928;
ROM1[1838]<=26'd1942813; ROM2[1838]<=26'd11288394; ROM3[1838]<=26'd9764123; ROM4[1838]<=26'd23467669;
ROM1[1839]<=26'd1942071; ROM2[1839]<=26'd11286629; ROM3[1839]<=26'd9761214; ROM4[1839]<=26'd23466254;
ROM1[1840]<=26'd1953459; ROM2[1840]<=26'd11288551; ROM3[1840]<=26'd9758099; ROM4[1840]<=26'd23467320;
ROM1[1841]<=26'd1969420; ROM2[1841]<=26'd11293125; ROM3[1841]<=26'd9754380; ROM4[1841]<=26'd23469153;
ROM1[1842]<=26'd1972106; ROM2[1842]<=26'd11292876; ROM3[1842]<=26'd9754258; ROM4[1842]<=26'd23468787;
ROM1[1843]<=26'd1962507; ROM2[1843]<=26'd11291229; ROM3[1843]<=26'd9754702; ROM4[1843]<=26'd23466834;
ROM1[1844]<=26'd1952600; ROM2[1844]<=26'd11289584; ROM3[1844]<=26'd9754312; ROM4[1844]<=26'd23464837;
ROM1[1845]<=26'd1945984; ROM2[1845]<=26'd11286073; ROM3[1845]<=26'd9756500; ROM4[1845]<=26'd23463571;
ROM1[1846]<=26'd1937899; ROM2[1846]<=26'd11284709; ROM3[1846]<=26'd9759701; ROM4[1846]<=26'd23463891;
ROM1[1847]<=26'd1939589; ROM2[1847]<=26'd11286021; ROM3[1847]<=26'd9762610; ROM4[1847]<=26'd23465424;
ROM1[1848]<=26'd1944357; ROM2[1848]<=26'd11283236; ROM3[1848]<=26'd9756820; ROM4[1848]<=26'd23462598;
ROM1[1849]<=26'd1955219; ROM2[1849]<=26'd11284562; ROM3[1849]<=26'd9750272; ROM4[1849]<=26'd23461315;
ROM1[1850]<=26'd1965019; ROM2[1850]<=26'd11287378; ROM3[1850]<=26'd9748621; ROM4[1850]<=26'd23462534;
ROM1[1851]<=26'd1958387; ROM2[1851]<=26'd11285930; ROM3[1851]<=26'd9748658; ROM4[1851]<=26'd23461675;
ROM1[1852]<=26'd1947845; ROM2[1852]<=26'd11282943; ROM3[1852]<=26'd9752542; ROM4[1852]<=26'd23462318;
ROM1[1853]<=26'd1947171; ROM2[1853]<=26'd11286780; ROM3[1853]<=26'd9759733; ROM4[1853]<=26'd23466006;
ROM1[1854]<=26'd1945345; ROM2[1854]<=26'd11291161; ROM3[1854]<=26'd9764637; ROM4[1854]<=26'd23469902;
ROM1[1855]<=26'd1942486; ROM2[1855]<=26'd11291972; ROM3[1855]<=26'd9766540; ROM4[1855]<=26'd23470024;
ROM1[1856]<=26'd1950633; ROM2[1856]<=26'd11295660; ROM3[1856]<=26'd9769128; ROM4[1856]<=26'd23471430;
ROM1[1857]<=26'd1962679; ROM2[1857]<=26'd11296795; ROM3[1857]<=26'd9765954; ROM4[1857]<=26'd23470635;
ROM1[1858]<=26'd1971314; ROM2[1858]<=26'd11296290; ROM3[1858]<=26'd9763477; ROM4[1858]<=26'd23469190;
ROM1[1859]<=26'd1972873; ROM2[1859]<=26'd11297791; ROM3[1859]<=26'd9765212; ROM4[1859]<=26'd23471352;
ROM1[1860]<=26'd1964375; ROM2[1860]<=26'd11296325; ROM3[1860]<=26'd9766795; ROM4[1860]<=26'd23470958;
ROM1[1861]<=26'd1956345; ROM2[1861]<=26'd11296367; ROM3[1861]<=26'd9769656; ROM4[1861]<=26'd23471173;
ROM1[1862]<=26'd1945649; ROM2[1862]<=26'd11289212; ROM3[1862]<=26'd9764775; ROM4[1862]<=26'd23465542;
ROM1[1863]<=26'd1933366; ROM2[1863]<=26'd11279924; ROM3[1863]<=26'd9760167; ROM4[1863]<=26'd23457867;
ROM1[1864]<=26'd1935215; ROM2[1864]<=26'd11280305; ROM3[1864]<=26'd9759392; ROM4[1864]<=26'd23456584;
ROM1[1865]<=26'd1947196; ROM2[1865]<=26'd11283828; ROM3[1865]<=26'd9756721; ROM4[1865]<=26'd23458451;
ROM1[1866]<=26'd1962466; ROM2[1866]<=26'd11286234; ROM3[1866]<=26'd9753275; ROM4[1866]<=26'd23459682;
ROM1[1867]<=26'd1961406; ROM2[1867]<=26'd11283493; ROM3[1867]<=26'd9748241; ROM4[1867]<=26'd23455519;
ROM1[1868]<=26'd1955618; ROM2[1868]<=26'd11283745; ROM3[1868]<=26'd9750811; ROM4[1868]<=26'd23457258;
ROM1[1869]<=26'd1952977; ROM2[1869]<=26'd11285829; ROM3[1869]<=26'd9760438; ROM4[1869]<=26'd23464366;
ROM1[1870]<=26'd1942235; ROM2[1870]<=26'd11280684; ROM3[1870]<=26'd9759404; ROM4[1870]<=26'd23461077;
ROM1[1871]<=26'd1940122; ROM2[1871]<=26'd11284419; ROM3[1871]<=26'd9766815; ROM4[1871]<=26'd23464871;
ROM1[1872]<=26'd1943820; ROM2[1872]<=26'd11288003; ROM3[1872]<=26'd9771887; ROM4[1872]<=26'd23468994;
ROM1[1873]<=26'd1933868; ROM2[1873]<=26'd11274332; ROM3[1873]<=26'd9753466; ROM4[1873]<=26'd23452408;
ROM1[1874]<=26'd1943451; ROM2[1874]<=26'd11273145; ROM3[1874]<=26'd9745903; ROM4[1874]<=26'd23448583;
ROM1[1875]<=26'd1951968; ROM2[1875]<=26'd11273953; ROM3[1875]<=26'd9743497; ROM4[1875]<=26'd23451460;
ROM1[1876]<=26'd1942559; ROM2[1876]<=26'd11268531; ROM3[1876]<=26'd9740263; ROM4[1876]<=26'd23446983;
ROM1[1877]<=26'd1936447; ROM2[1877]<=26'd11269061; ROM3[1877]<=26'd9745292; ROM4[1877]<=26'd23448374;
ROM1[1878]<=26'd1934269; ROM2[1878]<=26'd11273084; ROM3[1878]<=26'd9751304; ROM4[1878]<=26'd23452121;
ROM1[1879]<=26'd1929197; ROM2[1879]<=26'd11274791; ROM3[1879]<=26'd9757045; ROM4[1879]<=26'd23453877;
ROM1[1880]<=26'd1926149; ROM2[1880]<=26'd11274269; ROM3[1880]<=26'd9757463; ROM4[1880]<=26'd23453157;
ROM1[1881]<=26'd1932443; ROM2[1881]<=26'd11276125; ROM3[1881]<=26'd9755981; ROM4[1881]<=26'd23453000;
ROM1[1882]<=26'd1943998; ROM2[1882]<=26'd11278644; ROM3[1882]<=26'd9752396; ROM4[1882]<=26'd23452860;
ROM1[1883]<=26'd1954747; ROM2[1883]<=26'd11280921; ROM3[1883]<=26'd9747883; ROM4[1883]<=26'd23453800;
ROM1[1884]<=26'd1950404; ROM2[1884]<=26'd11277898; ROM3[1884]<=26'd9747082; ROM4[1884]<=26'd23453400;
ROM1[1885]<=26'd1943289; ROM2[1885]<=26'd11277059; ROM3[1885]<=26'd9752227; ROM4[1885]<=26'd23453926;
ROM1[1886]<=26'd1935901; ROM2[1886]<=26'd11273853; ROM3[1886]<=26'd9754252; ROM4[1886]<=26'd23452611;
ROM1[1887]<=26'd1929873; ROM2[1887]<=26'd11270550; ROM3[1887]<=26'd9755970; ROM4[1887]<=26'd23452315;
ROM1[1888]<=26'd1928811; ROM2[1888]<=26'd11275129; ROM3[1888]<=26'd9760657; ROM4[1888]<=26'd23456291;
ROM1[1889]<=26'd1932344; ROM2[1889]<=26'd11276925; ROM3[1889]<=26'd9759776; ROM4[1889]<=26'd23457322;
ROM1[1890]<=26'd1944124; ROM2[1890]<=26'd11279785; ROM3[1890]<=26'd9755859; ROM4[1890]<=26'd23457142;
ROM1[1891]<=26'd1960706; ROM2[1891]<=26'd11287284; ROM3[1891]<=26'd9755528; ROM4[1891]<=26'd23462384;
ROM1[1892]<=26'd1963162; ROM2[1892]<=26'd11285341; ROM3[1892]<=26'd9753969; ROM4[1892]<=26'd23462474;
ROM1[1893]<=26'd1957087; ROM2[1893]<=26'd11283599; ROM3[1893]<=26'd9755011; ROM4[1893]<=26'd23462810;
ROM1[1894]<=26'd1954704; ROM2[1894]<=26'd11288167; ROM3[1894]<=26'd9762700; ROM4[1894]<=26'd23469199;
ROM1[1895]<=26'd1951829; ROM2[1895]<=26'd11291003; ROM3[1895]<=26'd9766867; ROM4[1895]<=26'd23469961;
ROM1[1896]<=26'd1945378; ROM2[1896]<=26'd11289934; ROM3[1896]<=26'd9769172; ROM4[1896]<=26'd23468432;
ROM1[1897]<=26'd1949606; ROM2[1897]<=26'd11292426; ROM3[1897]<=26'd9773595; ROM4[1897]<=26'd23472331;
ROM1[1898]<=26'd1955449; ROM2[1898]<=26'd11293144; ROM3[1898]<=26'd9771563; ROM4[1898]<=26'd23471627;
ROM1[1899]<=26'd1963203; ROM2[1899]<=26'd11289648; ROM3[1899]<=26'd9762077; ROM4[1899]<=26'd23466864;
ROM1[1900]<=26'd1972164; ROM2[1900]<=26'd11294181; ROM3[1900]<=26'd9759807; ROM4[1900]<=26'd23469462;
ROM1[1901]<=26'd1965546; ROM2[1901]<=26'd11291393; ROM3[1901]<=26'd9756711; ROM4[1901]<=26'd23466662;
ROM1[1902]<=26'd1955118; ROM2[1902]<=26'd11286049; ROM3[1902]<=26'd9757057; ROM4[1902]<=26'd23463213;
ROM1[1903]<=26'd1950733; ROM2[1903]<=26'd11287090; ROM3[1903]<=26'd9760413; ROM4[1903]<=26'd23464379;
ROM1[1904]<=26'd1944849; ROM2[1904]<=26'd11286064; ROM3[1904]<=26'd9763000; ROM4[1904]<=26'd23464614;
ROM1[1905]<=26'd1941662; ROM2[1905]<=26'd11286867; ROM3[1905]<=26'd9766035; ROM4[1905]<=26'd23465106;
ROM1[1906]<=26'd1946878; ROM2[1906]<=26'd11287994; ROM3[1906]<=26'd9764536; ROM4[1906]<=26'd23464600;
ROM1[1907]<=26'd1957748; ROM2[1907]<=26'd11287629; ROM3[1907]<=26'd9758682; ROM4[1907]<=26'd23463576;
ROM1[1908]<=26'd1968835; ROM2[1908]<=26'd11289378; ROM3[1908]<=26'd9754885; ROM4[1908]<=26'd23463453;
ROM1[1909]<=26'd1967435; ROM2[1909]<=26'd11290768; ROM3[1909]<=26'd9755693; ROM4[1909]<=26'd23464456;
ROM1[1910]<=26'd1963032; ROM2[1910]<=26'd11293290; ROM3[1910]<=26'd9761210; ROM4[1910]<=26'd23469240;
ROM1[1911]<=26'd1960669; ROM2[1911]<=26'd11295825; ROM3[1911]<=26'd9767783; ROM4[1911]<=26'd23473245;
ROM1[1912]<=26'd1948049; ROM2[1912]<=26'd11291512; ROM3[1912]<=26'd9765836; ROM4[1912]<=26'd23467513;
ROM1[1913]<=26'd1941416; ROM2[1913]<=26'd11289938; ROM3[1913]<=26'd9766284; ROM4[1913]<=26'd23465254;
ROM1[1914]<=26'd1946368; ROM2[1914]<=26'd11293721; ROM3[1914]<=26'd9767716; ROM4[1914]<=26'd23467611;
ROM1[1915]<=26'd1959981; ROM2[1915]<=26'd11297907; ROM3[1915]<=26'd9766919; ROM4[1915]<=26'd23470629;
ROM1[1916]<=26'd1969726; ROM2[1916]<=26'd11294737; ROM3[1916]<=26'd9759123; ROM4[1916]<=26'd23465904;
ROM1[1917]<=26'd1962453; ROM2[1917]<=26'd11285037; ROM3[1917]<=26'd9749591; ROM4[1917]<=26'd23458111;
ROM1[1918]<=26'd1959148; ROM2[1918]<=26'd11288219; ROM3[1918]<=26'd9755790; ROM4[1918]<=26'd23462171;
ROM1[1919]<=26'd1953275; ROM2[1919]<=26'd11291774; ROM3[1919]<=26'd9763345; ROM4[1919]<=26'd23465403;
ROM1[1920]<=26'd1944459; ROM2[1920]<=26'd11288388; ROM3[1920]<=26'd9762017; ROM4[1920]<=26'd23463453;
ROM1[1921]<=26'd1941966; ROM2[1921]<=26'd11290579; ROM3[1921]<=26'd9767318; ROM4[1921]<=26'd23466410;
ROM1[1922]<=26'd1943246; ROM2[1922]<=26'd11290585; ROM3[1922]<=26'd9769863; ROM4[1922]<=26'd23468628;
ROM1[1923]<=26'd1946597; ROM2[1923]<=26'd11286485; ROM3[1923]<=26'd9764299; ROM4[1923]<=26'd23464718;
ROM1[1924]<=26'd1958904; ROM2[1924]<=26'd11287578; ROM3[1924]<=26'd9759203; ROM4[1924]<=26'd23464269;
ROM1[1925]<=26'd1969444; ROM2[1925]<=26'd11292004; ROM3[1925]<=26'd9758888; ROM4[1925]<=26'd23468116;
ROM1[1926]<=26'd1957967; ROM2[1926]<=26'd11284107; ROM3[1926]<=26'd9753027; ROM4[1926]<=26'd23461121;
ROM1[1927]<=26'd1943010; ROM2[1927]<=26'd11275549; ROM3[1927]<=26'd9746951; ROM4[1927]<=26'd23454403;
ROM1[1928]<=26'd1941425; ROM2[1928]<=26'd11279925; ROM3[1928]<=26'd9754831; ROM4[1928]<=26'd23459942;
ROM1[1929]<=26'd1933760; ROM2[1929]<=26'd11279523; ROM3[1929]<=26'd9758589; ROM4[1929]<=26'd23460718;
ROM1[1930]<=26'd1927599; ROM2[1930]<=26'd11277639; ROM3[1930]<=26'd9753813; ROM4[1930]<=26'd23456984;
ROM1[1931]<=26'd1931572; ROM2[1931]<=26'd11278541; ROM3[1931]<=26'd9750296; ROM4[1931]<=26'd23454141;
ROM1[1932]<=26'd1947345; ROM2[1932]<=26'd11280816; ROM3[1932]<=26'd9747088; ROM4[1932]<=26'd23454595;
ROM1[1933]<=26'd1961594; ROM2[1933]<=26'd11284481; ROM3[1933]<=26'd9745069; ROM4[1933]<=26'd23456552;
ROM1[1934]<=26'd1961585; ROM2[1934]<=26'd11286508; ROM3[1934]<=26'd9747347; ROM4[1934]<=26'd23458467;
ROM1[1935]<=26'd1956944; ROM2[1935]<=26'd11287970; ROM3[1935]<=26'd9753611; ROM4[1935]<=26'd23461512;
ROM1[1936]<=26'd1953308; ROM2[1936]<=26'd11290332; ROM3[1936]<=26'd9762388; ROM4[1936]<=26'd23465933;
ROM1[1937]<=26'd1953429; ROM2[1937]<=26'd11293680; ROM3[1937]<=26'd9769489; ROM4[1937]<=26'd23470970;
ROM1[1938]<=26'd1954309; ROM2[1938]<=26'd11298700; ROM3[1938]<=26'd9777703; ROM4[1938]<=26'd23477298;
ROM1[1939]<=26'd1953895; ROM2[1939]<=26'd11295452; ROM3[1939]<=26'd9775628; ROM4[1939]<=26'd23474760;
ROM1[1940]<=26'd1960560; ROM2[1940]<=26'd11291595; ROM3[1940]<=26'd9765927; ROM4[1940]<=26'd23470624;
ROM1[1941]<=26'd1970648; ROM2[1941]<=26'd11290092; ROM3[1941]<=26'd9757797; ROM4[1941]<=26'd23469125;
ROM1[1942]<=26'd1967187; ROM2[1942]<=26'd11285760; ROM3[1942]<=26'd9754400; ROM4[1942]<=26'd23466018;
ROM1[1943]<=26'd1962059; ROM2[1943]<=26'd11287047; ROM3[1943]<=26'd9760005; ROM4[1943]<=26'd23468012;
ROM1[1944]<=26'd1959337; ROM2[1944]<=26'd11290381; ROM3[1944]<=26'd9766418; ROM4[1944]<=26'd23470949;
ROM1[1945]<=26'd1957159; ROM2[1945]<=26'd11292398; ROM3[1945]<=26'd9772027; ROM4[1945]<=26'd23473965;
ROM1[1946]<=26'd1953228; ROM2[1946]<=26'd11292298; ROM3[1946]<=26'd9777756; ROM4[1946]<=26'd23476345;
ROM1[1947]<=26'd1951171; ROM2[1947]<=26'd11290874; ROM3[1947]<=26'd9777439; ROM4[1947]<=26'd23476442;
ROM1[1948]<=26'd1955629; ROM2[1948]<=26'd11287852; ROM3[1948]<=26'd9771264; ROM4[1948]<=26'd23474336;
ROM1[1949]<=26'd1964900; ROM2[1949]<=26'd11285391; ROM3[1949]<=26'd9762159; ROM4[1949]<=26'd23471433;
ROM1[1950]<=26'd1973018; ROM2[1950]<=26'd11286924; ROM3[1950]<=26'd9757469; ROM4[1950]<=26'd23469296;
ROM1[1951]<=26'd1970853; ROM2[1951]<=26'd11288554; ROM3[1951]<=26'd9758624; ROM4[1951]<=26'd23469067;
ROM1[1952]<=26'd1964347; ROM2[1952]<=26'd11291521; ROM3[1952]<=26'd9765038; ROM4[1952]<=26'd23472363;
ROM1[1953]<=26'd1964585; ROM2[1953]<=26'd11297696; ROM3[1953]<=26'd9773418; ROM4[1953]<=26'd23476313;
ROM1[1954]<=26'd1961495; ROM2[1954]<=26'd11300526; ROM3[1954]<=26'd9779353; ROM4[1954]<=26'd23479259;
ROM1[1955]<=26'd1954847; ROM2[1955]<=26'd11295473; ROM3[1955]<=26'd9776086; ROM4[1955]<=26'd23476440;
ROM1[1956]<=26'd1950717; ROM2[1956]<=26'd11286847; ROM3[1956]<=26'd9765060; ROM4[1956]<=26'd23466883;
ROM1[1957]<=26'd1956933; ROM2[1957]<=26'd11284632; ROM3[1957]<=26'd9755974; ROM4[1957]<=26'd23463171;
ROM1[1958]<=26'd1961985; ROM2[1958]<=26'd11280398; ROM3[1958]<=26'd9745282; ROM4[1958]<=26'd23457334;
ROM1[1959]<=26'd1963863; ROM2[1959]<=26'd11283242; ROM3[1959]<=26'd9746751; ROM4[1959]<=26'd23459480;
ROM1[1960]<=26'd1966328; ROM2[1960]<=26'd11292956; ROM3[1960]<=26'd9758498; ROM4[1960]<=26'd23470037;
ROM1[1961]<=26'd1959199; ROM2[1961]<=26'd11290013; ROM3[1961]<=26'd9759783; ROM4[1961]<=26'd23468635;
ROM1[1962]<=26'd1948124; ROM2[1962]<=26'd11285112; ROM3[1962]<=26'd9757254; ROM4[1962]<=26'd23465170;
ROM1[1963]<=26'd1943229; ROM2[1963]<=26'd11286476; ROM3[1963]<=26'd9760465; ROM4[1963]<=26'd23465125;
ROM1[1964]<=26'd1947174; ROM2[1964]<=26'd11287226; ROM3[1964]<=26'd9761096; ROM4[1964]<=26'd23465511;
ROM1[1965]<=26'd1959968; ROM2[1965]<=26'd11292307; ROM3[1965]<=26'd9759089; ROM4[1965]<=26'd23468094;
ROM1[1966]<=26'd1971951; ROM2[1966]<=26'd11291260; ROM3[1966]<=26'd9752306; ROM4[1966]<=26'd23466293;
ROM1[1967]<=26'd1967430; ROM2[1967]<=26'd11283589; ROM3[1967]<=26'd9743791; ROM4[1967]<=26'd23459648;
ROM1[1968]<=26'd1956823; ROM2[1968]<=26'd11280592; ROM3[1968]<=26'd9743424; ROM4[1968]<=26'd23455841;
ROM1[1969]<=26'd1948481; ROM2[1969]<=26'd11277574; ROM3[1969]<=26'd9745813; ROM4[1969]<=26'd23454680;
ROM1[1970]<=26'd1948200; ROM2[1970]<=26'd11281163; ROM3[1970]<=26'd9750869; ROM4[1970]<=26'd23459061;
ROM1[1971]<=26'd1944496; ROM2[1971]<=26'd11283709; ROM3[1971]<=26'd9755614; ROM4[1971]<=26'd23461501;
ROM1[1972]<=26'd1937580; ROM2[1972]<=26'd11278281; ROM3[1972]<=26'd9749110; ROM4[1972]<=26'd23455687;
ROM1[1973]<=26'd1940456; ROM2[1973]<=26'd11275149; ROM3[1973]<=26'd9742696; ROM4[1973]<=26'd23452086;
ROM1[1974]<=26'd1953539; ROM2[1974]<=26'd11277101; ROM3[1974]<=26'd9740250; ROM4[1974]<=26'd23452864;
ROM1[1975]<=26'd1961190; ROM2[1975]<=26'd11280402; ROM3[1975]<=26'd9740085; ROM4[1975]<=26'd23456474;
ROM1[1976]<=26'd1956859; ROM2[1976]<=26'd11281469; ROM3[1976]<=26'd9741935; ROM4[1976]<=26'd23457047;
ROM1[1977]<=26'd1945508; ROM2[1977]<=26'd11279470; ROM3[1977]<=26'd9744182; ROM4[1977]<=26'd23452520;
ROM1[1978]<=26'd1943725; ROM2[1978]<=26'd11282077; ROM3[1978]<=26'd9750020; ROM4[1978]<=26'd23456419;
ROM1[1979]<=26'd1941278; ROM2[1979]<=26'd11284121; ROM3[1979]<=26'd9755234; ROM4[1979]<=26'd23460550;
ROM1[1980]<=26'd1932824; ROM2[1980]<=26'd11280581; ROM3[1980]<=26'd9751060; ROM4[1980]<=26'd23456802;
ROM1[1981]<=26'd1939473; ROM2[1981]<=26'd11282393; ROM3[1981]<=26'd9749676; ROM4[1981]<=26'd23457178;
ROM1[1982]<=26'd1957482; ROM2[1982]<=26'd11289566; ROM3[1982]<=26'd9752566; ROM4[1982]<=26'd23461383;
ROM1[1983]<=26'd1973906; ROM2[1983]<=26'd11297434; ROM3[1983]<=26'd9752669; ROM4[1983]<=26'd23465925;
ROM1[1984]<=26'd1971674; ROM2[1984]<=26'd11295785; ROM3[1984]<=26'd9753822; ROM4[1984]<=26'd23465855;
ROM1[1985]<=26'd1958379; ROM2[1985]<=26'd11286926; ROM3[1985]<=26'd9750516; ROM4[1985]<=26'd23460064;
ROM1[1986]<=26'd1947739; ROM2[1986]<=26'd11284336; ROM3[1986]<=26'd9750321; ROM4[1986]<=26'd23456810;
ROM1[1987]<=26'd1933820; ROM2[1987]<=26'd11275519; ROM3[1987]<=26'd9745628; ROM4[1987]<=26'd23447350;
ROM1[1988]<=26'd1933068; ROM2[1988]<=26'd11274832; ROM3[1988]<=26'd9747312; ROM4[1988]<=26'd23448438;
ROM1[1989]<=26'd1939320; ROM2[1989]<=26'd11278077; ROM3[1989]<=26'd9749226; ROM4[1989]<=26'd23452232;
ROM1[1990]<=26'd1944598; ROM2[1990]<=26'd11274559; ROM3[1990]<=26'd9740458; ROM4[1990]<=26'd23447413;
ROM1[1991]<=26'd1956850; ROM2[1991]<=26'd11276900; ROM3[1991]<=26'd9735702; ROM4[1991]<=26'd23447636;
ROM1[1992]<=26'd1959116; ROM2[1992]<=26'd11278366; ROM3[1992]<=26'd9736364; ROM4[1992]<=26'd23447512;
ROM1[1993]<=26'd1954489; ROM2[1993]<=26'd11280425; ROM3[1993]<=26'd9739880; ROM4[1993]<=26'd23450341;
ROM1[1994]<=26'd1947877; ROM2[1994]<=26'd11280722; ROM3[1994]<=26'd9745945; ROM4[1994]<=26'd23452620;
ROM1[1995]<=26'd1945720; ROM2[1995]<=26'd11282028; ROM3[1995]<=26'd9752406; ROM4[1995]<=26'd23455522;
ROM1[1996]<=26'd1950487; ROM2[1996]<=26'd11290354; ROM3[1996]<=26'd9763614; ROM4[1996]<=26'd23465163;
ROM1[1997]<=26'd1948372; ROM2[1997]<=26'd11288303; ROM3[1997]<=26'd9763987; ROM4[1997]<=26'd23463917;
ROM1[1998]<=26'd1946324; ROM2[1998]<=26'd11278286; ROM3[1998]<=26'd9750547; ROM4[1998]<=26'd23452712;
ROM1[1999]<=26'd1960312; ROM2[1999]<=26'd11280022; ROM3[1999]<=26'd9744345; ROM4[1999]<=26'd23453159;
ROM1[2000]<=26'd1968851; ROM2[2000]<=26'd11286411; ROM3[2000]<=26'd9746693; ROM4[2000]<=26'd23459486;
ROM1[2001]<=26'd1966749; ROM2[2001]<=26'd11289111; ROM3[2001]<=26'd9751728; ROM4[2001]<=26'd23461411;
ROM1[2002]<=26'd1957487; ROM2[2002]<=26'd11284946; ROM3[2002]<=26'd9751440; ROM4[2002]<=26'd23458739;
ROM1[2003]<=26'd1948090; ROM2[2003]<=26'd11281986; ROM3[2003]<=26'd9751529; ROM4[2003]<=26'd23457223;
ROM1[2004]<=26'd1935860; ROM2[2004]<=26'd11274476; ROM3[2004]<=26'd9747791; ROM4[2004]<=26'd23449897;
ROM1[2005]<=26'd1930202; ROM2[2005]<=26'd11271293; ROM3[2005]<=26'd9744337; ROM4[2005]<=26'd23445408;
ROM1[2006]<=26'd1939907; ROM2[2006]<=26'd11277491; ROM3[2006]<=26'd9747661; ROM4[2006]<=26'd23451653;
ROM1[2007]<=26'd1955577; ROM2[2007]<=26'd11280925; ROM3[2007]<=26'd9746555; ROM4[2007]<=26'd23455011;
ROM1[2008]<=26'd1966550; ROM2[2008]<=26'd11282503; ROM3[2008]<=26'd9743244; ROM4[2008]<=26'd23456266;
ROM1[2009]<=26'd1962629; ROM2[2009]<=26'd11281862; ROM3[2009]<=26'd9744608; ROM4[2009]<=26'd23457624;
ROM1[2010]<=26'd1952933; ROM2[2010]<=26'd11280142; ROM3[2010]<=26'd9745687; ROM4[2010]<=26'd23455405;
ROM1[2011]<=26'd1941834; ROM2[2011]<=26'd11276533; ROM3[2011]<=26'd9744590; ROM4[2011]<=26'd23451717;
ROM1[2012]<=26'd1933464; ROM2[2012]<=26'd11272646; ROM3[2012]<=26'd9744806; ROM4[2012]<=26'd23450485;
ROM1[2013]<=26'd1929963; ROM2[2013]<=26'd11271586; ROM3[2013]<=26'd9748532; ROM4[2013]<=26'd23453851;
ROM1[2014]<=26'd1934173; ROM2[2014]<=26'd11274246; ROM3[2014]<=26'd9751033; ROM4[2014]<=26'd23457342;
ROM1[2015]<=26'd1945139; ROM2[2015]<=26'd11276352; ROM3[2015]<=26'd9749047; ROM4[2015]<=26'd23458279;
ROM1[2016]<=26'd1959218; ROM2[2016]<=26'd11278099; ROM3[2016]<=26'd9744266; ROM4[2016]<=26'd23458287;
ROM1[2017]<=26'd1962134; ROM2[2017]<=26'd11279329; ROM3[2017]<=26'd9743933; ROM4[2017]<=26'd23458816;
ROM1[2018]<=26'd1956991; ROM2[2018]<=26'd11279582; ROM3[2018]<=26'd9747871; ROM4[2018]<=26'd23460313;
ROM1[2019]<=26'd1950352; ROM2[2019]<=26'd11277393; ROM3[2019]<=26'd9750848; ROM4[2019]<=26'd23460368;
ROM1[2020]<=26'd1943430; ROM2[2020]<=26'd11275356; ROM3[2020]<=26'd9751758; ROM4[2020]<=26'd23458181;
ROM1[2021]<=26'd1937124; ROM2[2021]<=26'd11275792; ROM3[2021]<=26'd9753672; ROM4[2021]<=26'd23457055;
ROM1[2022]<=26'd1938802; ROM2[2022]<=26'd11278761; ROM3[2022]<=26'd9753735; ROM4[2022]<=26'd23458796;
ROM1[2023]<=26'd1946887; ROM2[2023]<=26'd11281071; ROM3[2023]<=26'd9751533; ROM4[2023]<=26'd23458573;
ROM1[2024]<=26'd1961218; ROM2[2024]<=26'd11282294; ROM3[2024]<=26'd9748464; ROM4[2024]<=26'd23459288;
ROM1[2025]<=26'd1966620; ROM2[2025]<=26'd11280909; ROM3[2025]<=26'd9743410; ROM4[2025]<=26'd23457842;
ROM1[2026]<=26'd1958805; ROM2[2026]<=26'd11278143; ROM3[2026]<=26'd9741546; ROM4[2026]<=26'd23455203;
ROM1[2027]<=26'd1953694; ROM2[2027]<=26'd11281144; ROM3[2027]<=26'd9747049; ROM4[2027]<=26'd23457941;
ROM1[2028]<=26'd1955092; ROM2[2028]<=26'd11287174; ROM3[2028]<=26'd9757799; ROM4[2028]<=26'd23465393;
ROM1[2029]<=26'd1955801; ROM2[2029]<=26'd11293241; ROM3[2029]<=26'd9766873; ROM4[2029]<=26'd23471624;
ROM1[2030]<=26'd1948132; ROM2[2030]<=26'd11289433; ROM3[2030]<=26'd9763989; ROM4[2030]<=26'd23468160;
ROM1[2031]<=26'd1948108; ROM2[2031]<=26'd11283610; ROM3[2031]<=26'd9758837; ROM4[2031]<=26'd23464517;
ROM1[2032]<=26'd1960719; ROM2[2032]<=26'd11285008; ROM3[2032]<=26'd9754824; ROM4[2032]<=26'd23463854;
ROM1[2033]<=26'd1969229; ROM2[2033]<=26'd11283646; ROM3[2033]<=26'd9746554; ROM4[2033]<=26'd23461616;
ROM1[2034]<=26'd1969030; ROM2[2034]<=26'd11285487; ROM3[2034]<=26'd9749848; ROM4[2034]<=26'd23464067;
ROM1[2035]<=26'd1965865; ROM2[2035]<=26'd11289175; ROM3[2035]<=26'd9756232; ROM4[2035]<=26'd23467984;
ROM1[2036]<=26'd1959902; ROM2[2036]<=26'd11291559; ROM3[2036]<=26'd9758881; ROM4[2036]<=26'd23469728;
ROM1[2037]<=26'd1955154; ROM2[2037]<=26'd11292529; ROM3[2037]<=26'd9763394; ROM4[2037]<=26'd23470667;
ROM1[2038]<=26'd1948011; ROM2[2038]<=26'd11287401; ROM3[2038]<=26'd9760136; ROM4[2038]<=26'd23466795;
ROM1[2039]<=26'd1943073; ROM2[2039]<=26'd11278173; ROM3[2039]<=26'd9751178; ROM4[2039]<=26'd23457545;
ROM1[2040]<=26'd1947275; ROM2[2040]<=26'd11272282; ROM3[2040]<=26'd9742329; ROM4[2040]<=26'd23449917;
ROM1[2041]<=26'd1961393; ROM2[2041]<=26'd11278233; ROM3[2041]<=26'd9740667; ROM4[2041]<=26'd23453739;
ROM1[2042]<=26'd1977289; ROM2[2042]<=26'd11291516; ROM3[2042]<=26'd9754277; ROM4[2042]<=26'd23467310;
ROM1[2043]<=26'd1972041; ROM2[2043]<=26'd11291594; ROM3[2043]<=26'd9758517; ROM4[2043]<=26'd23468994;
ROM1[2044]<=26'd1951050; ROM2[2044]<=26'd11278421; ROM3[2044]<=26'd9749357; ROM4[2044]<=26'd23457763;
ROM1[2045]<=26'd1938949; ROM2[2045]<=26'd11272280; ROM3[2045]<=26'd9745727; ROM4[2045]<=26'd23451427;
ROM1[2046]<=26'd1929019; ROM2[2046]<=26'd11268329; ROM3[2046]<=26'd9746338; ROM4[2046]<=26'd23447774;
ROM1[2047]<=26'd1929686; ROM2[2047]<=26'd11270792; ROM3[2047]<=26'd9748376; ROM4[2047]<=26'd23449379;
ROM1[2048]<=26'd1944418; ROM2[2048]<=26'd11278644; ROM3[2048]<=26'd9750021; ROM4[2048]<=26'd23454520;
ROM1[2049]<=26'd1961418; ROM2[2049]<=26'd11282722; ROM3[2049]<=26'd9746466; ROM4[2049]<=26'd23455830;
ROM1[2050]<=26'd1963203; ROM2[2050]<=26'd11280386; ROM3[2050]<=26'd9738623; ROM4[2050]<=26'd23451213;
ROM1[2051]<=26'd1957769; ROM2[2051]<=26'd11279176; ROM3[2051]<=26'd9739370; ROM4[2051]<=26'd23450464;
ROM1[2052]<=26'd1952640; ROM2[2052]<=26'd11281152; ROM3[2052]<=26'd9744577; ROM4[2052]<=26'd23453152;
ROM1[2053]<=26'd1947261; ROM2[2053]<=26'd11280467; ROM3[2053]<=26'd9748650; ROM4[2053]<=26'd23454002;
ROM1[2054]<=26'd1941309; ROM2[2054]<=26'd11278674; ROM3[2054]<=26'd9751101; ROM4[2054]<=26'd23453698;
ROM1[2055]<=26'd1939732; ROM2[2055]<=26'd11279843; ROM3[2055]<=26'd9751233; ROM4[2055]<=26'd23453041;
ROM1[2056]<=26'd1947546; ROM2[2056]<=26'd11284226; ROM3[2056]<=26'd9752154; ROM4[2056]<=26'd23456390;
ROM1[2057]<=26'd1959300; ROM2[2057]<=26'd11285515; ROM3[2057]<=26'd9745610; ROM4[2057]<=26'd23455853;
ROM1[2058]<=26'd1966919; ROM2[2058]<=26'd11282954; ROM3[2058]<=26'd9736883; ROM4[2058]<=26'd23452336;
ROM1[2059]<=26'd1965447; ROM2[2059]<=26'd11283076; ROM3[2059]<=26'd9737459; ROM4[2059]<=26'd23453416;
ROM1[2060]<=26'd1959602; ROM2[2060]<=26'd11284697; ROM3[2060]<=26'd9740658; ROM4[2060]<=26'd23454569;
ROM1[2061]<=26'd1956070; ROM2[2061]<=26'd11286485; ROM3[2061]<=26'd9747756; ROM4[2061]<=26'd23458141;
ROM1[2062]<=26'd1955373; ROM2[2062]<=26'd11290424; ROM3[2062]<=26'd9755626; ROM4[2062]<=26'd23464033;
ROM1[2063]<=26'd1945224; ROM2[2063]<=26'd11285243; ROM3[2063]<=26'd9753447; ROM4[2063]<=26'd23460169;
ROM1[2064]<=26'd1943545; ROM2[2064]<=26'd11282187; ROM3[2064]<=26'd9749364; ROM4[2064]<=26'd23457305;
ROM1[2065]<=26'd1951949; ROM2[2065]<=26'd11282452; ROM3[2065]<=26'd9743835; ROM4[2065]<=26'd23454384;
ROM1[2066]<=26'd1966511; ROM2[2066]<=26'd11287051; ROM3[2066]<=26'd9742515; ROM4[2066]<=26'd23457109;
ROM1[2067]<=26'd1970747; ROM2[2067]<=26'd11290703; ROM3[2067]<=26'd9744464; ROM4[2067]<=26'd23461379;
ROM1[2068]<=26'd1961123; ROM2[2068]<=26'd11286952; ROM3[2068]<=26'd9743442; ROM4[2068]<=26'd23459466;
ROM1[2069]<=26'd1953832; ROM2[2069]<=26'd11287370; ROM3[2069]<=26'd9746345; ROM4[2069]<=26'd23460023;
ROM1[2070]<=26'd1948998; ROM2[2070]<=26'd11287768; ROM3[2070]<=26'd9748484; ROM4[2070]<=26'd23459677;
ROM1[2071]<=26'd1945992; ROM2[2071]<=26'd11289253; ROM3[2071]<=26'd9752238; ROM4[2071]<=26'd23460298;
ROM1[2072]<=26'd1945830; ROM2[2072]<=26'd11287023; ROM3[2072]<=26'd9751254; ROM4[2072]<=26'd23457720;
ROM1[2073]<=26'd1952718; ROM2[2073]<=26'd11285827; ROM3[2073]<=26'd9747432; ROM4[2073]<=26'd23457205;
ROM1[2074]<=26'd1962799; ROM2[2074]<=26'd11288367; ROM3[2074]<=26'd9741312; ROM4[2074]<=26'd23456402;
ROM1[2075]<=26'd1967492; ROM2[2075]<=26'd11288175; ROM3[2075]<=26'd9738333; ROM4[2075]<=26'd23456555;
ROM1[2076]<=26'd1964023; ROM2[2076]<=26'd11287457; ROM3[2076]<=26'd9743353; ROM4[2076]<=26'd23458569;
ROM1[2077]<=26'd1952388; ROM2[2077]<=26'd11283856; ROM3[2077]<=26'd9743668; ROM4[2077]<=26'd23454493;
ROM1[2078]<=26'd1944774; ROM2[2078]<=26'd11279959; ROM3[2078]<=26'd9745644; ROM4[2078]<=26'd23453693;
ROM1[2079]<=26'd1938580; ROM2[2079]<=26'd11278922; ROM3[2079]<=26'd9746999; ROM4[2079]<=26'd23453525;
ROM1[2080]<=26'd1937018; ROM2[2080]<=26'd11280242; ROM3[2080]<=26'd9748655; ROM4[2080]<=26'd23455454;
ROM1[2081]<=26'd1943275; ROM2[2081]<=26'd11281370; ROM3[2081]<=26'd9750310; ROM4[2081]<=26'd23458291;
ROM1[2082]<=26'd1954284; ROM2[2082]<=26'd11281975; ROM3[2082]<=26'd9744933; ROM4[2082]<=26'd23456195;
ROM1[2083]<=26'd1962991; ROM2[2083]<=26'd11279825; ROM3[2083]<=26'd9741435; ROM4[2083]<=26'd23455984;
ROM1[2084]<=26'd1960714; ROM2[2084]<=26'd11281103; ROM3[2084]<=26'd9744390; ROM4[2084]<=26'd23458601;
ROM1[2085]<=26'd1954018; ROM2[2085]<=26'd11281145; ROM3[2085]<=26'd9748209; ROM4[2085]<=26'd23459830;
ROM1[2086]<=26'd1955087; ROM2[2086]<=26'd11285556; ROM3[2086]<=26'd9757271; ROM4[2086]<=26'd23464875;
ROM1[2087]<=26'd1961417; ROM2[2087]<=26'd11298724; ROM3[2087]<=26'd9772269; ROM4[2087]<=26'd23478040;
ROM1[2088]<=26'd1961011; ROM2[2088]<=26'd11304541; ROM3[2088]<=26'd9778785; ROM4[2088]<=26'd23482474;
ROM1[2089]<=26'd1953275; ROM2[2089]<=26'd11294850; ROM3[2089]<=26'd9767654; ROM4[2089]<=26'd23471577;
ROM1[2090]<=26'd1949787; ROM2[2090]<=26'd11283979; ROM3[2090]<=26'd9750190; ROM4[2090]<=26'd23458858;
ROM1[2091]<=26'd1952153; ROM2[2091]<=26'd11277133; ROM3[2091]<=26'd9733407; ROM4[2091]<=26'd23448349;
ROM1[2092]<=26'd1947127; ROM2[2092]<=26'd11269458; ROM3[2092]<=26'd9726288; ROM4[2092]<=26'd23442014;
ROM1[2093]<=26'd1947738; ROM2[2093]<=26'd11275452; ROM3[2093]<=26'd9736362; ROM4[2093]<=26'd23449659;
ROM1[2094]<=26'd1945912; ROM2[2094]<=26'd11280103; ROM3[2094]<=26'd9747220; ROM4[2094]<=26'd23457461;
ROM1[2095]<=26'd1938951; ROM2[2095]<=26'd11276783; ROM3[2095]<=26'd9750367; ROM4[2095]<=26'd23457173;
ROM1[2096]<=26'd1931754; ROM2[2096]<=26'd11274329; ROM3[2096]<=26'd9750371; ROM4[2096]<=26'd23453986;
ROM1[2097]<=26'd1931972; ROM2[2097]<=26'd11273516; ROM3[2097]<=26'd9748475; ROM4[2097]<=26'd23451496;
ROM1[2098]<=26'd1942459; ROM2[2098]<=26'd11274018; ROM3[2098]<=26'd9746517; ROM4[2098]<=26'd23451800;
ROM1[2099]<=26'd1958959; ROM2[2099]<=26'd11279743; ROM3[2099]<=26'd9743705; ROM4[2099]<=26'd23454700;
ROM1[2100]<=26'd1968632; ROM2[2100]<=26'd11285596; ROM3[2100]<=26'd9744460; ROM4[2100]<=26'd23458663;
ROM1[2101]<=26'd1962811; ROM2[2101]<=26'd11284506; ROM3[2101]<=26'd9746797; ROM4[2101]<=26'd23461211;
ROM1[2102]<=26'd1952602; ROM2[2102]<=26'd11279987; ROM3[2102]<=26'd9745605; ROM4[2102]<=26'd23458789;
ROM1[2103]<=26'd1949000; ROM2[2103]<=26'd11280560; ROM3[2103]<=26'd9751008; ROM4[2103]<=26'd23459449;
ROM1[2104]<=26'd1951012; ROM2[2104]<=26'd11288265; ROM3[2104]<=26'd9762228; ROM4[2104]<=26'd23467646;
ROM1[2105]<=26'd1946432; ROM2[2105]<=26'd11285582; ROM3[2105]<=26'd9761512; ROM4[2105]<=26'd23463725;
ROM1[2106]<=26'd1947514; ROM2[2106]<=26'd11283771; ROM3[2106]<=26'd9758459; ROM4[2106]<=26'd23460949;
ROM1[2107]<=26'd1960293; ROM2[2107]<=26'd11287042; ROM3[2107]<=26'd9753423; ROM4[2107]<=26'd23460589;
ROM1[2108]<=26'd1963974; ROM2[2108]<=26'd11282161; ROM3[2108]<=26'd9741617; ROM4[2108]<=26'd23453328;
ROM1[2109]<=26'd1962991; ROM2[2109]<=26'd11283117; ROM3[2109]<=26'd9742883; ROM4[2109]<=26'd23455118;
ROM1[2110]<=26'd1960064; ROM2[2110]<=26'd11285914; ROM3[2110]<=26'd9750732; ROM4[2110]<=26'd23459277;
ROM1[2111]<=26'd1949895; ROM2[2111]<=26'd11281188; ROM3[2111]<=26'd9750980; ROM4[2111]<=26'd23455922;
ROM1[2112]<=26'd1946948; ROM2[2112]<=26'd11283436; ROM3[2112]<=26'd9755430; ROM4[2112]<=26'd23459140;
ROM1[2113]<=26'd1949095; ROM2[2113]<=26'd11288647; ROM3[2113]<=26'd9762571; ROM4[2113]<=26'd23465781;
ROM1[2114]<=26'd1947500; ROM2[2114]<=26'd11285489; ROM3[2114]<=26'd9755510; ROM4[2114]<=26'd23460952;
ROM1[2115]<=26'd1950405; ROM2[2115]<=26'd11279693; ROM3[2115]<=26'd9742253; ROM4[2115]<=26'd23453422;
ROM1[2116]<=26'd1962601; ROM2[2116]<=26'd11279651; ROM3[2116]<=26'd9738428; ROM4[2116]<=26'd23453662;
ROM1[2117]<=26'd1959675; ROM2[2117]<=26'd11278420; ROM3[2117]<=26'd9735260; ROM4[2117]<=26'd23451962;
ROM1[2118]<=26'd1950788; ROM2[2118]<=26'd11276309; ROM3[2118]<=26'd9735224; ROM4[2118]<=26'd23451551;
ROM1[2119]<=26'd1950833; ROM2[2119]<=26'd11281555; ROM3[2119]<=26'd9746153; ROM4[2119]<=26'd23459085;
ROM1[2120]<=26'd1943646; ROM2[2120]<=26'd11278631; ROM3[2120]<=26'd9747149; ROM4[2120]<=26'd23458222;
ROM1[2121]<=26'd1933951; ROM2[2121]<=26'd11273173; ROM3[2121]<=26'd9745557; ROM4[2121]<=26'd23453640;
ROM1[2122]<=26'd1940353; ROM2[2122]<=26'd11280276; ROM3[2122]<=26'd9752735; ROM4[2122]<=26'd23461354;
ROM1[2123]<=26'd1946759; ROM2[2123]<=26'd11280620; ROM3[2123]<=26'd9749125; ROM4[2123]<=26'd23461183;
ROM1[2124]<=26'd1952246; ROM2[2124]<=26'd11272864; ROM3[2124]<=26'd9734539; ROM4[2124]<=26'd23452941;
ROM1[2125]<=26'd1959046; ROM2[2125]<=26'd11274736; ROM3[2125]<=26'd9731293; ROM4[2125]<=26'd23454324;
ROM1[2126]<=26'd1954632; ROM2[2126]<=26'd11274470; ROM3[2126]<=26'd9734342; ROM4[2126]<=26'd23454022;
ROM1[2127]<=26'd1948002; ROM2[2127]<=26'd11273477; ROM3[2127]<=26'd9738697; ROM4[2127]<=26'd23454925;
ROM1[2128]<=26'd1946459; ROM2[2128]<=26'd11278343; ROM3[2128]<=26'd9745938; ROM4[2128]<=26'd23459768;
ROM1[2129]<=26'd1945911; ROM2[2129]<=26'd11280657; ROM3[2129]<=26'd9753202; ROM4[2129]<=26'd23464768;
ROM1[2130]<=26'd1947006; ROM2[2130]<=26'd11282036; ROM3[2130]<=26'd9756555; ROM4[2130]<=26'd23468181;
ROM1[2131]<=26'd1952693; ROM2[2131]<=26'd11284186; ROM3[2131]<=26'd9756157; ROM4[2131]<=26'd23469011;
ROM1[2132]<=26'd1963354; ROM2[2132]<=26'd11284943; ROM3[2132]<=26'd9751883; ROM4[2132]<=26'd23468008;
ROM1[2133]<=26'd1970667; ROM2[2133]<=26'd11285946; ROM3[2133]<=26'd9744906; ROM4[2133]<=26'd23466154;
ROM1[2134]<=26'd1965725; ROM2[2134]<=26'd11285682; ROM3[2134]<=26'd9744282; ROM4[2134]<=26'd23464079;
ROM1[2135]<=26'd1958208; ROM2[2135]<=26'd11284820; ROM3[2135]<=26'd9748679; ROM4[2135]<=26'd23462616;
ROM1[2136]<=26'd1954252; ROM2[2136]<=26'd11287757; ROM3[2136]<=26'd9755163; ROM4[2136]<=26'd23465282;
ROM1[2137]<=26'd1950682; ROM2[2137]<=26'd11286709; ROM3[2137]<=26'd9759968; ROM4[2137]<=26'd23466462;
ROM1[2138]<=26'd1947683; ROM2[2138]<=26'd11283873; ROM3[2138]<=26'd9762211; ROM4[2138]<=26'd23464944;
ROM1[2139]<=26'd1947002; ROM2[2139]<=26'd11281090; ROM3[2139]<=26'd9759206; ROM4[2139]<=26'd23463909;
ROM1[2140]<=26'd1956765; ROM2[2140]<=26'd11282972; ROM3[2140]<=26'd9756535; ROM4[2140]<=26'd23464213;
ROM1[2141]<=26'd1971680; ROM2[2141]<=26'd11289852; ROM3[2141]<=26'd9756643; ROM4[2141]<=26'd23468493;
ROM1[2142]<=26'd1969021; ROM2[2142]<=26'd11288232; ROM3[2142]<=26'd9753069; ROM4[2142]<=26'd23466147;
ROM1[2143]<=26'd1958732; ROM2[2143]<=26'd11284483; ROM3[2143]<=26'd9752275; ROM4[2143]<=26'd23463102;
ROM1[2144]<=26'd1951205; ROM2[2144]<=26'd11282321; ROM3[2144]<=26'd9755650; ROM4[2144]<=26'd23462560;
ROM1[2145]<=26'd1944561; ROM2[2145]<=26'd11278511; ROM3[2145]<=26'd9755239; ROM4[2145]<=26'd23459801;
ROM1[2146]<=26'd1942643; ROM2[2146]<=26'd11281229; ROM3[2146]<=26'd9758326; ROM4[2146]<=26'd23462672;
ROM1[2147]<=26'd1946736; ROM2[2147]<=26'd11284500; ROM3[2147]<=26'd9759771; ROM4[2147]<=26'd23464437;
ROM1[2148]<=26'd1949742; ROM2[2148]<=26'd11280022; ROM3[2148]<=26'd9750275; ROM4[2148]<=26'd23459429;
ROM1[2149]<=26'd1961816; ROM2[2149]<=26'd11281492; ROM3[2149]<=26'd9745253; ROM4[2149]<=26'd23459550;
ROM1[2150]<=26'd1971556; ROM2[2150]<=26'd11286798; ROM3[2150]<=26'd9748551; ROM4[2150]<=26'd23464456;
ROM1[2151]<=26'd1966180; ROM2[2151]<=26'd11287124; ROM3[2151]<=26'd9751862; ROM4[2151]<=26'd23465301;
ROM1[2152]<=26'd1964600; ROM2[2152]<=26'd11290123; ROM3[2152]<=26'd9758974; ROM4[2152]<=26'd23469278;
ROM1[2153]<=26'd1956366; ROM2[2153]<=26'd11283653; ROM3[2153]<=26'd9758088; ROM4[2153]<=26'd23464681;
ROM1[2154]<=26'd1944748; ROM2[2154]<=26'd11278658; ROM3[2154]<=26'd9758891; ROM4[2154]<=26'd23462973;
ROM1[2155]<=26'd1948407; ROM2[2155]<=26'd11283153; ROM3[2155]<=26'd9767995; ROM4[2155]<=26'd23471299;
ROM1[2156]<=26'd1952932; ROM2[2156]<=26'd11282242; ROM3[2156]<=26'd9765884; ROM4[2156]<=26'd23470315;
ROM1[2157]<=26'd1964489; ROM2[2157]<=26'd11283068; ROM3[2157]<=26'd9758669; ROM4[2157]<=26'd23468451;
ROM1[2158]<=26'd1978085; ROM2[2158]<=26'd11286191; ROM3[2158]<=26'd9755340; ROM4[2158]<=26'd23470746;
ROM1[2159]<=26'd1969676; ROM2[2159]<=26'd11280580; ROM3[2159]<=26'd9749551; ROM4[2159]<=26'd23464890;
ROM1[2160]<=26'd1957694; ROM2[2160]<=26'd11276100; ROM3[2160]<=26'd9749530; ROM4[2160]<=26'd23462269;
ROM1[2161]<=26'd1957533; ROM2[2161]<=26'd11280962; ROM3[2161]<=26'd9759864; ROM4[2161]<=26'd23468747;
ROM1[2162]<=26'd1949184; ROM2[2162]<=26'd11277340; ROM3[2162]<=26'd9757437; ROM4[2162]<=26'd23465613;
ROM1[2163]<=26'd1934990; ROM2[2163]<=26'd11267809; ROM3[2163]<=26'd9748569; ROM4[2163]<=26'd23455648;
ROM1[2164]<=26'd1936137; ROM2[2164]<=26'd11267824; ROM3[2164]<=26'd9748592; ROM4[2164]<=26'd23454901;
ROM1[2165]<=26'd1945792; ROM2[2165]<=26'd11268482; ROM3[2165]<=26'd9743410; ROM4[2165]<=26'd23454344;
ROM1[2166]<=26'd1957111; ROM2[2166]<=26'd11267652; ROM3[2166]<=26'd9737832; ROM4[2166]<=26'd23452303;
ROM1[2167]<=26'd1961230; ROM2[2167]<=26'd11270782; ROM3[2167]<=26'd9740371; ROM4[2167]<=26'd23455116;
ROM1[2168]<=26'd1957405; ROM2[2168]<=26'd11272751; ROM3[2168]<=26'd9742714; ROM4[2168]<=26'd23457305;
ROM1[2169]<=26'd1950735; ROM2[2169]<=26'd11272383; ROM3[2169]<=26'd9745415; ROM4[2169]<=26'd23457536;
ROM1[2170]<=26'd1946388; ROM2[2170]<=26'd11274338; ROM3[2170]<=26'd9749056; ROM4[2170]<=26'd23457784;
ROM1[2171]<=26'd1947303; ROM2[2171]<=26'd11278794; ROM3[2171]<=26'd9755507; ROM4[2171]<=26'd23464082;
ROM1[2172]<=26'd1949057; ROM2[2172]<=26'd11279776; ROM3[2172]<=26'd9756808; ROM4[2172]<=26'd23465787;
ROM1[2173]<=26'd1953174; ROM2[2173]<=26'd11278788; ROM3[2173]<=26'd9752197; ROM4[2173]<=26'd23462466;
ROM1[2174]<=26'd1967685; ROM2[2174]<=26'd11281250; ROM3[2174]<=26'd9748245; ROM4[2174]<=26'd23463718;
ROM1[2175]<=26'd1976167; ROM2[2175]<=26'd11283150; ROM3[2175]<=26'd9746656; ROM4[2175]<=26'd23465902;
ROM1[2176]<=26'd1965389; ROM2[2176]<=26'd11278046; ROM3[2176]<=26'd9742573; ROM4[2176]<=26'd23462011;
ROM1[2177]<=26'd1956725; ROM2[2177]<=26'd11277858; ROM3[2177]<=26'd9745581; ROM4[2177]<=26'd23463176;
ROM1[2178]<=26'd1957494; ROM2[2178]<=26'd11284730; ROM3[2178]<=26'd9754385; ROM4[2178]<=26'd23469153;
ROM1[2179]<=26'd1949473; ROM2[2179]<=26'd11283768; ROM3[2179]<=26'd9754911; ROM4[2179]<=26'd23466387;
ROM1[2180]<=26'd1950303; ROM2[2180]<=26'd11285812; ROM3[2180]<=26'd9758237; ROM4[2180]<=26'd23469128;
ROM1[2181]<=26'd1962180; ROM2[2181]<=26'd11290341; ROM3[2181]<=26'd9760144; ROM4[2181]<=26'd23473107;
ROM1[2182]<=26'd1965811; ROM2[2182]<=26'd11280842; ROM3[2182]<=26'd9747154; ROM4[2182]<=26'd23463765;
ROM1[2183]<=26'd1970907; ROM2[2183]<=26'd11277642; ROM3[2183]<=26'd9740705; ROM4[2183]<=26'd23460122;
ROM1[2184]<=26'd1968288; ROM2[2184]<=26'd11278554; ROM3[2184]<=26'd9742242; ROM4[2184]<=26'd23460978;
ROM1[2185]<=26'd1958569; ROM2[2185]<=26'd11274940; ROM3[2185]<=26'd9742435; ROM4[2185]<=26'd23459856;
ROM1[2186]<=26'd1954354; ROM2[2186]<=26'd11276043; ROM3[2186]<=26'd9746608; ROM4[2186]<=26'd23461903;
ROM1[2187]<=26'd1953719; ROM2[2187]<=26'd11279299; ROM3[2187]<=26'd9752620; ROM4[2187]<=26'd23465528;
ROM1[2188]<=26'd1951393; ROM2[2188]<=26'd11280747; ROM3[2188]<=26'd9755750; ROM4[2188]<=26'd23466818;
ROM1[2189]<=26'd1948805; ROM2[2189]<=26'd11277578; ROM3[2189]<=26'd9750568; ROM4[2189]<=26'd23461317;
ROM1[2190]<=26'd1956237; ROM2[2190]<=26'd11277541; ROM3[2190]<=26'd9744092; ROM4[2190]<=26'd23458208;
ROM1[2191]<=26'd1968290; ROM2[2191]<=26'd11280060; ROM3[2191]<=26'd9739222; ROM4[2191]<=26'd23458512;
ROM1[2192]<=26'd1970224; ROM2[2192]<=26'd11279462; ROM3[2192]<=26'd9736900; ROM4[2192]<=26'd23458389;
ROM1[2193]<=26'd1964146; ROM2[2193]<=26'd11279845; ROM3[2193]<=26'd9740438; ROM4[2193]<=26'd23461326;
ROM1[2194]<=26'd1955179; ROM2[2194]<=26'd11278089; ROM3[2194]<=26'd9744199; ROM4[2194]<=26'd23461736;
ROM1[2195]<=26'd1947621; ROM2[2195]<=26'd11274256; ROM3[2195]<=26'd9745755; ROM4[2195]<=26'd23458600;
ROM1[2196]<=26'd1942392; ROM2[2196]<=26'd11273640; ROM3[2196]<=26'd9747785; ROM4[2196]<=26'd23457191;
ROM1[2197]<=26'd1943076; ROM2[2197]<=26'd11273445; ROM3[2197]<=26'd9748769; ROM4[2197]<=26'd23456961;
ROM1[2198]<=26'd1951271; ROM2[2198]<=26'd11276490; ROM3[2198]<=26'd9749203; ROM4[2198]<=26'd23458517;
ROM1[2199]<=26'd1964894; ROM2[2199]<=26'd11278156; ROM3[2199]<=26'd9742974; ROM4[2199]<=26'd23458777;
ROM1[2200]<=26'd1970176; ROM2[2200]<=26'd11277763; ROM3[2200]<=26'd9740682; ROM4[2200]<=26'd23457187;
ROM1[2201]<=26'd1963325; ROM2[2201]<=26'd11276883; ROM3[2201]<=26'd9742694; ROM4[2201]<=26'd23455977;
ROM1[2202]<=26'd1957574; ROM2[2202]<=26'd11278314; ROM3[2202]<=26'd9746592; ROM4[2202]<=26'd23458592;
ROM1[2203]<=26'd1957404; ROM2[2203]<=26'd11281335; ROM3[2203]<=26'd9753548; ROM4[2203]<=26'd23462964;
ROM1[2204]<=26'd1947586; ROM2[2204]<=26'd11277563; ROM3[2204]<=26'd9751998; ROM4[2204]<=26'd23460789;
ROM1[2205]<=26'd1940517; ROM2[2205]<=26'd11273568; ROM3[2205]<=26'd9749077; ROM4[2205]<=26'd23456607;
ROM1[2206]<=26'd1946390; ROM2[2206]<=26'd11273352; ROM3[2206]<=26'd9745451; ROM4[2206]<=26'd23455261;
ROM1[2207]<=26'd1957251; ROM2[2207]<=26'd11274321; ROM3[2207]<=26'd9738369; ROM4[2207]<=26'd23454156;
ROM1[2208]<=26'd1963759; ROM2[2208]<=26'd11274240; ROM3[2208]<=26'd9734430; ROM4[2208]<=26'd23451762;
ROM1[2209]<=26'd1961738; ROM2[2209]<=26'd11275472; ROM3[2209]<=26'd9735748; ROM4[2209]<=26'd23453209;
ROM1[2210]<=26'd1950291; ROM2[2210]<=26'd11271727; ROM3[2210]<=26'd9734491; ROM4[2210]<=26'd23451383;
ROM1[2211]<=26'd1942117; ROM2[2211]<=26'd11270932; ROM3[2211]<=26'd9738632; ROM4[2211]<=26'd23452470;
ROM1[2212]<=26'd1938617; ROM2[2212]<=26'd11272628; ROM3[2212]<=26'd9742672; ROM4[2212]<=26'd23455146;
ROM1[2213]<=26'd1928668; ROM2[2213]<=26'd11264442; ROM3[2213]<=26'd9736107; ROM4[2213]<=26'd23447790;
ROM1[2214]<=26'd1927682; ROM2[2214]<=26'd11260532; ROM3[2214]<=26'd9732380; ROM4[2214]<=26'd23443232;
ROM1[2215]<=26'd1939807; ROM2[2215]<=26'd11262140; ROM3[2215]<=26'd9730875; ROM4[2215]<=26'd23444237;
ROM1[2216]<=26'd1955552; ROM2[2216]<=26'd11267794; ROM3[2216]<=26'd9732275; ROM4[2216]<=26'd23450357;
ROM1[2217]<=26'd1963266; ROM2[2217]<=26'd11276428; ROM3[2217]<=26'd9740251; ROM4[2217]<=26'd23459407;
ROM1[2218]<=26'd1962003; ROM2[2218]<=26'd11280781; ROM3[2218]<=26'd9748399; ROM4[2218]<=26'd23464767;
ROM1[2219]<=26'd1954289; ROM2[2219]<=26'd11279933; ROM3[2219]<=26'd9752833; ROM4[2219]<=26'd23464599;
ROM1[2220]<=26'd1943281; ROM2[2220]<=26'd11274211; ROM3[2220]<=26'd9749973; ROM4[2220]<=26'd23458032;
ROM1[2221]<=26'd1934566; ROM2[2221]<=26'd11270654; ROM3[2221]<=26'd9749590; ROM4[2221]<=26'd23454968;
ROM1[2222]<=26'd1936574; ROM2[2222]<=26'd11271395; ROM3[2222]<=26'd9750403; ROM4[2222]<=26'd23457047;
ROM1[2223]<=26'd1943880; ROM2[2223]<=26'd11273187; ROM3[2223]<=26'd9745186; ROM4[2223]<=26'd23455832;
ROM1[2224]<=26'd1956360; ROM2[2224]<=26'd11273973; ROM3[2224]<=26'd9738169; ROM4[2224]<=26'd23455949;
ROM1[2225]<=26'd1965050; ROM2[2225]<=26'd11276363; ROM3[2225]<=26'd9737721; ROM4[2225]<=26'd23458955;
ROM1[2226]<=26'd1961312; ROM2[2226]<=26'd11279381; ROM3[2226]<=26'd9741109; ROM4[2226]<=26'd23461121;
ROM1[2227]<=26'd1952673; ROM2[2227]<=26'd11278665; ROM3[2227]<=26'd9742337; ROM4[2227]<=26'd23461653;
ROM1[2228]<=26'd1949740; ROM2[2228]<=26'd11279077; ROM3[2228]<=26'd9744287; ROM4[2228]<=26'd23462098;
ROM1[2229]<=26'd1944508; ROM2[2229]<=26'd11278506; ROM3[2229]<=26'd9746146; ROM4[2229]<=26'd23460992;
ROM1[2230]<=26'd1939162; ROM2[2230]<=26'd11276205; ROM3[2230]<=26'd9744035; ROM4[2230]<=26'd23457579;
ROM1[2231]<=26'd1942394; ROM2[2231]<=26'd11275600; ROM3[2231]<=26'd9740967; ROM4[2231]<=26'd23454901;
ROM1[2232]<=26'd1952592; ROM2[2232]<=26'd11277371; ROM3[2232]<=26'd9738192; ROM4[2232]<=26'd23454048;
ROM1[2233]<=26'd1961951; ROM2[2233]<=26'd11279027; ROM3[2233]<=26'd9735365; ROM4[2233]<=26'd23454768;
ROM1[2234]<=26'd1959350; ROM2[2234]<=26'd11277491; ROM3[2234]<=26'd9736751; ROM4[2234]<=26'd23452959;
ROM1[2235]<=26'd1947420; ROM2[2235]<=26'd11272081; ROM3[2235]<=26'd9733752; ROM4[2235]<=26'd23447258;
ROM1[2236]<=26'd1940958; ROM2[2236]<=26'd11270395; ROM3[2236]<=26'd9734441; ROM4[2236]<=26'd23445888;
ROM1[2237]<=26'd1934356; ROM2[2237]<=26'd11270083; ROM3[2237]<=26'd9735102; ROM4[2237]<=26'd23444378;
ROM1[2238]<=26'd1928372; ROM2[2238]<=26'd11269738; ROM3[2238]<=26'd9733712; ROM4[2238]<=26'd23443327;
ROM1[2239]<=26'd1933543; ROM2[2239]<=26'd11271315; ROM3[2239]<=26'd9735564; ROM4[2239]<=26'd23446032;
ROM1[2240]<=26'd1942272; ROM2[2240]<=26'd11271184; ROM3[2240]<=26'd9731164; ROM4[2240]<=26'd23445779;
ROM1[2241]<=26'd1954522; ROM2[2241]<=26'd11273403; ROM3[2241]<=26'd9725565; ROM4[2241]<=26'd23445363;
ROM1[2242]<=26'd1963239; ROM2[2242]<=26'd11279913; ROM3[2242]<=26'd9730341; ROM4[2242]<=26'd23452179;
ROM1[2243]<=26'd1959491; ROM2[2243]<=26'd11282035; ROM3[2243]<=26'd9733685; ROM4[2243]<=26'd23455571;
ROM1[2244]<=26'd1947394; ROM2[2244]<=26'd11275715; ROM3[2244]<=26'd9732015; ROM4[2244]<=26'd23450709;
ROM1[2245]<=26'd1940776; ROM2[2245]<=26'd11273073; ROM3[2245]<=26'd9734869; ROM4[2245]<=26'd23450160;
ROM1[2246]<=26'd1930883; ROM2[2246]<=26'd11267566; ROM3[2246]<=26'd9732036; ROM4[2246]<=26'd23445828;
ROM1[2247]<=26'd1928381; ROM2[2247]<=26'd11265634; ROM3[2247]<=26'd9730669; ROM4[2247]<=26'd23443770;
ROM1[2248]<=26'd1940915; ROM2[2248]<=26'd11271758; ROM3[2248]<=26'd9732716; ROM4[2248]<=26'd23448710;
ROM1[2249]<=26'd1953025; ROM2[2249]<=26'd11270863; ROM3[2249]<=26'd9724780; ROM4[2249]<=26'd23447235;
ROM1[2250]<=26'd1951760; ROM2[2250]<=26'd11264383; ROM3[2250]<=26'd9716729; ROM4[2250]<=26'd23441542;
ROM1[2251]<=26'd1948517; ROM2[2251]<=26'd11266326; ROM3[2251]<=26'd9720943; ROM4[2251]<=26'd23443030;
ROM1[2252]<=26'd1949361; ROM2[2252]<=26'd11272728; ROM3[2252]<=26'd9731810; ROM4[2252]<=26'd23450726;
ROM1[2253]<=26'd1941474; ROM2[2253]<=26'd11269806; ROM3[2253]<=26'd9732362; ROM4[2253]<=26'd23448344;
ROM1[2254]<=26'd1930154; ROM2[2254]<=26'd11263606; ROM3[2254]<=26'd9730623; ROM4[2254]<=26'd23444203;
ROM1[2255]<=26'd1928389; ROM2[2255]<=26'd11263140; ROM3[2255]<=26'd9732471; ROM4[2255]<=26'd23444680;
ROM1[2256]<=26'd1932716; ROM2[2256]<=26'd11263232; ROM3[2256]<=26'd9728364; ROM4[2256]<=26'd23441653;
ROM1[2257]<=26'd1945407; ROM2[2257]<=26'd11266106; ROM3[2257]<=26'd9724067; ROM4[2257]<=26'd23442217;
ROM1[2258]<=26'd1955869; ROM2[2258]<=26'd11270710; ROM3[2258]<=26'd9722104; ROM4[2258]<=26'd23445570;
ROM1[2259]<=26'd1953057; ROM2[2259]<=26'd11269883; ROM3[2259]<=26'd9724030; ROM4[2259]<=26'd23446648;
ROM1[2260]<=26'd1942090; ROM2[2260]<=26'd11263293; ROM3[2260]<=26'd9725168; ROM4[2260]<=26'd23443417;
ROM1[2261]<=26'd1932078; ROM2[2261]<=26'd11260137; ROM3[2261]<=26'd9724846; ROM4[2261]<=26'd23440536;
ROM1[2262]<=26'd1930120; ROM2[2262]<=26'd11264335; ROM3[2262]<=26'd9730517; ROM4[2262]<=26'd23443630;
ROM1[2263]<=26'd1930957; ROM2[2263]<=26'd11268121; ROM3[2263]<=26'd9734830; ROM4[2263]<=26'd23446032;
ROM1[2264]<=26'd1938687; ROM2[2264]<=26'd11276190; ROM3[2264]<=26'd9738591; ROM4[2264]<=26'd23452048;
ROM1[2265]<=26'd1950223; ROM2[2265]<=26'd11279331; ROM3[2265]<=26'd9737131; ROM4[2265]<=26'd23454755;
ROM1[2266]<=26'd1953477; ROM2[2266]<=26'd11269323; ROM3[2266]<=26'd9723823; ROM4[2266]<=26'd23445699;
ROM1[2267]<=26'd1947286; ROM2[2267]<=26'd11263099; ROM3[2267]<=26'd9715755; ROM4[2267]<=26'd23438299;
ROM1[2268]<=26'd1938122; ROM2[2268]<=26'd11261010; ROM3[2268]<=26'd9714587; ROM4[2268]<=26'd23435546;
ROM1[2269]<=26'd1931978; ROM2[2269]<=26'd11261969; ROM3[2269]<=26'd9721213; ROM4[2269]<=26'd23437768;
ROM1[2270]<=26'd1930955; ROM2[2270]<=26'd11268569; ROM3[2270]<=26'd9729855; ROM4[2270]<=26'd23442798;
ROM1[2271]<=26'd1927323; ROM2[2271]<=26'd11271013; ROM3[2271]<=26'd9736460; ROM4[2271]<=26'd23446464;
ROM1[2272]<=26'd1925715; ROM2[2272]<=26'd11268950; ROM3[2272]<=26'd9733405; ROM4[2272]<=26'd23443794;
ROM1[2273]<=26'd1928767; ROM2[2273]<=26'd11265262; ROM3[2273]<=26'd9721672; ROM4[2273]<=26'd23435405;
ROM1[2274]<=26'd1942868; ROM2[2274]<=26'd11267893; ROM3[2274]<=26'd9716123; ROM4[2274]<=26'd23434569;
ROM1[2275]<=26'd1944457; ROM2[2275]<=26'd11265335; ROM3[2275]<=26'd9709470; ROM4[2275]<=26'd23431883;
ROM1[2276]<=26'd1936778; ROM2[2276]<=26'd11263035; ROM3[2276]<=26'd9712091; ROM4[2276]<=26'd23431406;
ROM1[2277]<=26'd1936564; ROM2[2277]<=26'd11270857; ROM3[2277]<=26'd9725918; ROM4[2277]<=26'd23441007;
ROM1[2278]<=26'd1936088; ROM2[2278]<=26'd11276817; ROM3[2278]<=26'd9734962; ROM4[2278]<=26'd23447776;
ROM1[2279]<=26'd1937535; ROM2[2279]<=26'd11283341; ROM3[2279]<=26'd9743104; ROM4[2279]<=26'd23454461;
ROM1[2280]<=26'd1936647; ROM2[2280]<=26'd11283922; ROM3[2280]<=26'd9743346; ROM4[2280]<=26'd23454517;
ROM1[2281]<=26'd1934596; ROM2[2281]<=26'd11276503; ROM3[2281]<=26'd9734146; ROM4[2281]<=26'd23447846;
ROM1[2282]<=26'd1938054; ROM2[2282]<=26'd11267625; ROM3[2282]<=26'd9721024; ROM4[2282]<=26'd23438378;
ROM1[2283]<=26'd1941329; ROM2[2283]<=26'd11262407; ROM3[2283]<=26'd9713544; ROM4[2283]<=26'd23433651;
ROM1[2284]<=26'd1939133; ROM2[2284]<=26'd11262031; ROM3[2284]<=26'd9716472; ROM4[2284]<=26'd23434849;
ROM1[2285]<=26'd1934935; ROM2[2285]<=26'd11263440; ROM3[2285]<=26'd9722805; ROM4[2285]<=26'd23436545;
ROM1[2286]<=26'd1931418; ROM2[2286]<=26'd11264606; ROM3[2286]<=26'd9728952; ROM4[2286]<=26'd23438887;
ROM1[2287]<=26'd1923223; ROM2[2287]<=26'd11263078; ROM3[2287]<=26'd9730668; ROM4[2287]<=26'd23437563;
ROM1[2288]<=26'd1915985; ROM2[2288]<=26'd11261257; ROM3[2288]<=26'd9730202; ROM4[2288]<=26'd23435563;
ROM1[2289]<=26'd1916916; ROM2[2289]<=26'd11260273; ROM3[2289]<=26'd9728912; ROM4[2289]<=26'd23434495;
ROM1[2290]<=26'd1931506; ROM2[2290]<=26'd11266765; ROM3[2290]<=26'd9727964; ROM4[2290]<=26'd23438421;
ROM1[2291]<=26'd1950817; ROM2[2291]<=26'd11276719; ROM3[2291]<=26'd9726975; ROM4[2291]<=26'd23443851;
ROM1[2292]<=26'd1947220; ROM2[2292]<=26'd11273700; ROM3[2292]<=26'd9723018; ROM4[2292]<=26'd23440505;
ROM1[2293]<=26'd1937259; ROM2[2293]<=26'd11268473; ROM3[2293]<=26'd9721171; ROM4[2293]<=26'd23436177;
ROM1[2294]<=26'd1929674; ROM2[2294]<=26'd11266000; ROM3[2294]<=26'd9725021; ROM4[2294]<=26'd23436179;
ROM1[2295]<=26'd1922344; ROM2[2295]<=26'd11262671; ROM3[2295]<=26'd9727437; ROM4[2295]<=26'd23435742;
ROM1[2296]<=26'd1921626; ROM2[2296]<=26'd11266381; ROM3[2296]<=26'd9733366; ROM4[2296]<=26'd23440478;
ROM1[2297]<=26'd1925946; ROM2[2297]<=26'd11270623; ROM3[2297]<=26'd9737568; ROM4[2297]<=26'd23445467;
ROM1[2298]<=26'd1933576; ROM2[2298]<=26'd11273078; ROM3[2298]<=26'd9734309; ROM4[2298]<=26'd23445539;
ROM1[2299]<=26'd1944869; ROM2[2299]<=26'd11272389; ROM3[2299]<=26'd9727291; ROM4[2299]<=26'd23443998;
ROM1[2300]<=26'd1945990; ROM2[2300]<=26'd11267089; ROM3[2300]<=26'd9720508; ROM4[2300]<=26'd23440122;
ROM1[2301]<=26'd1942177; ROM2[2301]<=26'd11268834; ROM3[2301]<=26'd9722891; ROM4[2301]<=26'd23443495;
ROM1[2302]<=26'd1940708; ROM2[2302]<=26'd11272671; ROM3[2302]<=26'd9731813; ROM4[2302]<=26'd23449259;
ROM1[2303]<=26'd1934491; ROM2[2303]<=26'd11270489; ROM3[2303]<=26'd9732953; ROM4[2303]<=26'd23447282;
ROM1[2304]<=26'd1929783; ROM2[2304]<=26'd11271921; ROM3[2304]<=26'd9736533; ROM4[2304]<=26'd23450099;
ROM1[2305]<=26'd1932264; ROM2[2305]<=26'd11275848; ROM3[2305]<=26'd9743121; ROM4[2305]<=26'd23454456;
ROM1[2306]<=26'd1932698; ROM2[2306]<=26'd11272077; ROM3[2306]<=26'd9737953; ROM4[2306]<=26'd23448930;
ROM1[2307]<=26'd1943746; ROM2[2307]<=26'd11271875; ROM3[2307]<=26'd9732284; ROM4[2307]<=26'd23448456;
ROM1[2308]<=26'd1955693; ROM2[2308]<=26'd11275200; ROM3[2308]<=26'd9730780; ROM4[2308]<=26'd23451221;
ROM1[2309]<=26'd1953005; ROM2[2309]<=26'd11273603; ROM3[2309]<=26'd9731624; ROM4[2309]<=26'd23450886;
ROM1[2310]<=26'd1949583; ROM2[2310]<=26'd11276304; ROM3[2310]<=26'd9736765; ROM4[2310]<=26'd23455106;
ROM1[2311]<=26'd1942302; ROM2[2311]<=26'd11275289; ROM3[2311]<=26'd9739476; ROM4[2311]<=26'd23453417;
ROM1[2312]<=26'd1935586; ROM2[2312]<=26'd11275121; ROM3[2312]<=26'd9741423; ROM4[2312]<=26'd23452947;
ROM1[2313]<=26'd1936410; ROM2[2313]<=26'd11281880; ROM3[2313]<=26'd9748593; ROM4[2313]<=26'd23458836;
ROM1[2314]<=26'd1939691; ROM2[2314]<=26'd11283680; ROM3[2314]<=26'd9749316; ROM4[2314]<=26'd23459883;
ROM1[2315]<=26'd1947935; ROM2[2315]<=26'd11283695; ROM3[2315]<=26'd9742602; ROM4[2315]<=26'd23458872;
ROM1[2316]<=26'd1955398; ROM2[2316]<=26'd11280472; ROM3[2316]<=26'd9734702; ROM4[2316]<=26'd23454059;
ROM1[2317]<=26'd1949526; ROM2[2317]<=26'd11274115; ROM3[2317]<=26'd9725687; ROM4[2317]<=26'd23445262;
ROM1[2318]<=26'd1934180; ROM2[2318]<=26'd11262914; ROM3[2318]<=26'd9719081; ROM4[2318]<=26'd23436182;
ROM1[2319]<=26'd1929312; ROM2[2319]<=26'd11262600; ROM3[2319]<=26'd9725148; ROM4[2319]<=26'd23437413;
ROM1[2320]<=26'd1937030; ROM2[2320]<=26'd11273742; ROM3[2320]<=26'd9735230; ROM4[2320]<=26'd23447611;
ROM1[2321]<=26'd1924101; ROM2[2321]<=26'd11266226; ROM3[2321]<=26'd9730365; ROM4[2321]<=26'd23441346;
ROM1[2322]<=26'd1916990; ROM2[2322]<=26'd11260411; ROM3[2322]<=26'd9725892; ROM4[2322]<=26'd23436565;
ROM1[2323]<=26'd1923523; ROM2[2323]<=26'd11259612; ROM3[2323]<=26'd9722434; ROM4[2323]<=26'd23435552;
ROM1[2324]<=26'd1935324; ROM2[2324]<=26'd11256694; ROM3[2324]<=26'd9716402; ROM4[2324]<=26'd23432840;
ROM1[2325]<=26'd1947464; ROM2[2325]<=26'd11263660; ROM3[2325]<=26'd9719008; ROM4[2325]<=26'd23438069;
ROM1[2326]<=26'd1946441; ROM2[2326]<=26'd11268499; ROM3[2326]<=26'd9722676; ROM4[2326]<=26'd23441683;
ROM1[2327]<=26'd1938913; ROM2[2327]<=26'd11267700; ROM3[2327]<=26'd9726939; ROM4[2327]<=26'd23442747;
ROM1[2328]<=26'd1931964; ROM2[2328]<=26'd11266736; ROM3[2328]<=26'd9731344; ROM4[2328]<=26'd23444022;
ROM1[2329]<=26'd1925895; ROM2[2329]<=26'd11266283; ROM3[2329]<=26'd9736130; ROM4[2329]<=26'd23444977;
ROM1[2330]<=26'd1923839; ROM2[2330]<=26'd11267565; ROM3[2330]<=26'd9736353; ROM4[2330]<=26'd23443951;
ROM1[2331]<=26'd1930026; ROM2[2331]<=26'd11268403; ROM3[2331]<=26'd9732791; ROM4[2331]<=26'd23443363;
ROM1[2332]<=26'd1940484; ROM2[2332]<=26'd11267192; ROM3[2332]<=26'd9725678; ROM4[2332]<=26'd23440050;
ROM1[2333]<=26'd1948007; ROM2[2333]<=26'd11266351; ROM3[2333]<=26'd9718179; ROM4[2333]<=26'd23437568;
ROM1[2334]<=26'd1948183; ROM2[2334]<=26'd11268238; ROM3[2334]<=26'd9721185; ROM4[2334]<=26'd23440296;
ROM1[2335]<=26'd1935320; ROM2[2335]<=26'd11263776; ROM3[2335]<=26'd9720092; ROM4[2335]<=26'd23436032;
ROM1[2336]<=26'd1927359; ROM2[2336]<=26'd11260616; ROM3[2336]<=26'd9721351; ROM4[2336]<=26'd23433296;
ROM1[2337]<=26'd1922915; ROM2[2337]<=26'd11259530; ROM3[2337]<=26'd9726738; ROM4[2337]<=26'd23434564;
ROM1[2338]<=26'd1922833; ROM2[2338]<=26'd11263382; ROM3[2338]<=26'd9734594; ROM4[2338]<=26'd23438837;
ROM1[2339]<=26'd1931550; ROM2[2339]<=26'd11268028; ROM3[2339]<=26'd9738419; ROM4[2339]<=26'd23444945;
ROM1[2340]<=26'd1933556; ROM2[2340]<=26'd11262114; ROM3[2340]<=26'd9727033; ROM4[2340]<=26'd23438200;
ROM1[2341]<=26'd1945321; ROM2[2341]<=26'd11263892; ROM3[2341]<=26'd9722133; ROM4[2341]<=26'd23437062;
ROM1[2342]<=26'd1949134; ROM2[2342]<=26'd11265013; ROM3[2342]<=26'd9723025; ROM4[2342]<=26'd23441229;
ROM1[2343]<=26'd1941753; ROM2[2343]<=26'd11263810; ROM3[2343]<=26'd9725389; ROM4[2343]<=26'd23441474;
ROM1[2344]<=26'd1939899; ROM2[2344]<=26'd11268313; ROM3[2344]<=26'd9734260; ROM4[2344]<=26'd23447299;
ROM1[2345]<=26'd1937051; ROM2[2345]<=26'd11269524; ROM3[2345]<=26'd9738860; ROM4[2345]<=26'd23450738;
ROM1[2346]<=26'd1929434; ROM2[2346]<=26'd11267037; ROM3[2346]<=26'd9740408; ROM4[2346]<=26'd23448922;
ROM1[2347]<=26'd1932349; ROM2[2347]<=26'd11271102; ROM3[2347]<=26'd9747142; ROM4[2347]<=26'd23451797;
ROM1[2348]<=26'd1942884; ROM2[2348]<=26'd11275651; ROM3[2348]<=26'd9746727; ROM4[2348]<=26'd23454327;
ROM1[2349]<=26'd1951003; ROM2[2349]<=26'd11270677; ROM3[2349]<=26'd9734972; ROM4[2349]<=26'd23450229;
ROM1[2350]<=26'd1951257; ROM2[2350]<=26'd11264342; ROM3[2350]<=26'd9728863; ROM4[2350]<=26'd23444396;
ROM1[2351]<=26'd1945424; ROM2[2351]<=26'd11261303; ROM3[2351]<=26'd9728977; ROM4[2351]<=26'd23441289;
ROM1[2352]<=26'd1938252; ROM2[2352]<=26'd11260353; ROM3[2352]<=26'd9732367; ROM4[2352]<=26'd23442316;
ROM1[2353]<=26'd1935464; ROM2[2353]<=26'd11263498; ROM3[2353]<=26'd9738131; ROM4[2353]<=26'd23446326;
ROM1[2354]<=26'd1929555; ROM2[2354]<=26'd11264881; ROM3[2354]<=26'd9741549; ROM4[2354]<=26'd23448491;
ROM1[2355]<=26'd1924783; ROM2[2355]<=26'd11264020; ROM3[2355]<=26'd9741124; ROM4[2355]<=26'd23447496;
ROM1[2356]<=26'd1932068; ROM2[2356]<=26'd11265789; ROM3[2356]<=26'd9740549; ROM4[2356]<=26'd23448878;
ROM1[2357]<=26'd1947686; ROM2[2357]<=26'd11270504; ROM3[2357]<=26'd9737985; ROM4[2357]<=26'd23450491;
ROM1[2358]<=26'd1961339; ROM2[2358]<=26'd11276095; ROM3[2358]<=26'd9737005; ROM4[2358]<=26'd23453843;
ROM1[2359]<=26'd1963504; ROM2[2359]<=26'd11280207; ROM3[2359]<=26'd9740072; ROM4[2359]<=26'd23458976;
ROM1[2360]<=26'd1952286; ROM2[2360]<=26'd11278044; ROM3[2360]<=26'd9739552; ROM4[2360]<=26'd23454643;
ROM1[2361]<=26'd1934944; ROM2[2361]<=26'd11267475; ROM3[2361]<=26'd9731046; ROM4[2361]<=26'd23443830;
ROM1[2362]<=26'd1925730; ROM2[2362]<=26'd11262536; ROM3[2362]<=26'd9725486; ROM4[2362]<=26'd23439243;
ROM1[2363]<=26'd1923318; ROM2[2363]<=26'd11266280; ROM3[2363]<=26'd9729683; ROM4[2363]<=26'd23442531;
ROM1[2364]<=26'd1930530; ROM2[2364]<=26'd11271487; ROM3[2364]<=26'd9734629; ROM4[2364]<=26'd23447426;
ROM1[2365]<=26'd1940173; ROM2[2365]<=26'd11271800; ROM3[2365]<=26'd9729730; ROM4[2365]<=26'd23446328;
ROM1[2366]<=26'd1949388; ROM2[2366]<=26'd11271708; ROM3[2366]<=26'd9723903; ROM4[2366]<=26'd23444392;
ROM1[2367]<=26'd1950017; ROM2[2367]<=26'd11270242; ROM3[2367]<=26'd9721224; ROM4[2367]<=26'd23442053;
ROM1[2368]<=26'd1944894; ROM2[2368]<=26'd11271941; ROM3[2368]<=26'd9726312; ROM4[2368]<=26'd23443944;
ROM1[2369]<=26'd1946756; ROM2[2369]<=26'd11280398; ROM3[2369]<=26'd9741749; ROM4[2369]<=26'd23454114;
ROM1[2370]<=26'd1944534; ROM2[2370]<=26'd11280505; ROM3[2370]<=26'd9747316; ROM4[2370]<=26'd23457854;
ROM1[2371]<=26'd1933434; ROM2[2371]<=26'd11276021; ROM3[2371]<=26'd9744314; ROM4[2371]<=26'd23453451;
ROM1[2372]<=26'd1932456; ROM2[2372]<=26'd11275969; ROM3[2372]<=26'd9741933; ROM4[2372]<=26'd23451418;
ROM1[2373]<=26'd1948387; ROM2[2373]<=26'd11283522; ROM3[2373]<=26'd9747109; ROM4[2373]<=26'd23459461;
ROM1[2374]<=26'd1966753; ROM2[2374]<=26'd11289764; ROM3[2374]<=26'd9750030; ROM4[2374]<=26'd23465433;
ROM1[2375]<=26'd1966685; ROM2[2375]<=26'd11284738; ROM3[2375]<=26'd9745212; ROM4[2375]<=26'd23460616;
ROM1[2376]<=26'd1949835; ROM2[2376]<=26'd11271357; ROM3[2376]<=26'd9735030; ROM4[2376]<=26'd23450192;
ROM1[2377]<=26'd1937227; ROM2[2377]<=26'd11267886; ROM3[2377]<=26'd9732217; ROM4[2377]<=26'd23447128;
ROM1[2378]<=26'd1935808; ROM2[2378]<=26'd11273921; ROM3[2378]<=26'd9739515; ROM4[2378]<=26'd23451646;
ROM1[2379]<=26'd1935739; ROM2[2379]<=26'd11278351; ROM3[2379]<=26'd9748464; ROM4[2379]<=26'd23457229;
ROM1[2380]<=26'd1942512; ROM2[2380]<=26'd11287093; ROM3[2380]<=26'd9758647; ROM4[2380]<=26'd23467500;
ROM1[2381]<=26'd1944405; ROM2[2381]<=26'd11284182; ROM3[2381]<=26'd9753389; ROM4[2381]<=26'd23463943;
ROM1[2382]<=26'd1948739; ROM2[2382]<=26'd11277505; ROM3[2382]<=26'd9741672; ROM4[2382]<=26'd23455656;
ROM1[2383]<=26'd1958349; ROM2[2383]<=26'd11279435; ROM3[2383]<=26'd9737481; ROM4[2383]<=26'd23457920;
ROM1[2384]<=26'd1956723; ROM2[2384]<=26'd11280189; ROM3[2384]<=26'd9736683; ROM4[2384]<=26'd23457214;
ROM1[2385]<=26'd1950037; ROM2[2385]<=26'd11279418; ROM3[2385]<=26'd9739262; ROM4[2385]<=26'd23455551;
ROM1[2386]<=26'd1947609; ROM2[2386]<=26'd11280313; ROM3[2386]<=26'd9744461; ROM4[2386]<=26'd23457421;
ROM1[2387]<=26'd1943361; ROM2[2387]<=26'd11279555; ROM3[2387]<=26'd9747398; ROM4[2387]<=26'd23457758;
ROM1[2388]<=26'd1936251; ROM2[2388]<=26'd11275280; ROM3[2388]<=26'd9746225; ROM4[2388]<=26'd23454731;
ROM1[2389]<=26'd1939198; ROM2[2389]<=26'd11274901; ROM3[2389]<=26'd9745346; ROM4[2389]<=26'd23454640;
ROM1[2390]<=26'd1948175; ROM2[2390]<=26'd11272685; ROM3[2390]<=26'd9737934; ROM4[2390]<=26'd23451802;
ROM1[2391]<=26'd1959650; ROM2[2391]<=26'd11273419; ROM3[2391]<=26'd9731093; ROM4[2391]<=26'd23449085;
ROM1[2392]<=26'd1962509; ROM2[2392]<=26'd11277789; ROM3[2392]<=26'd9737213; ROM4[2392]<=26'd23453626;
ROM1[2393]<=26'd1957402; ROM2[2393]<=26'd11280454; ROM3[2393]<=26'd9743656; ROM4[2393]<=26'd23457094;
ROM1[2394]<=26'd1945234; ROM2[2394]<=26'd11276373; ROM3[2394]<=26'd9742365; ROM4[2394]<=26'd23453861;
ROM1[2395]<=26'd1933659; ROM2[2395]<=26'd11269808; ROM3[2395]<=26'd9740044; ROM4[2395]<=26'd23450137;
ROM1[2396]<=26'd1926917; ROM2[2396]<=26'd11266630; ROM3[2396]<=26'd9739191; ROM4[2396]<=26'd23447866;
ROM1[2397]<=26'd1926024; ROM2[2397]<=26'd11265107; ROM3[2397]<=26'd9736114; ROM4[2397]<=26'd23444781;
ROM1[2398]<=26'd1934370; ROM2[2398]<=26'd11267461; ROM3[2398]<=26'd9733334; ROM4[2398]<=26'd23444030;
ROM1[2399]<=26'd1948757; ROM2[2399]<=26'd11269778; ROM3[2399]<=26'd9729103; ROM4[2399]<=26'd23445381;
ROM1[2400]<=26'd1953694; ROM2[2400]<=26'd11270035; ROM3[2400]<=26'd9728239; ROM4[2400]<=26'd23445506;
ROM1[2401]<=26'd1950880; ROM2[2401]<=26'd11270368; ROM3[2401]<=26'd9732887; ROM4[2401]<=26'd23447458;
ROM1[2402]<=26'd1943070; ROM2[2402]<=26'd11269458; ROM3[2402]<=26'd9737350; ROM4[2402]<=26'd23448288;
ROM1[2403]<=26'd1938355; ROM2[2403]<=26'd11270990; ROM3[2403]<=26'd9742406; ROM4[2403]<=26'd23449471;
ROM1[2404]<=26'd1938094; ROM2[2404]<=26'd11274995; ROM3[2404]<=26'd9749349; ROM4[2404]<=26'd23455328;
ROM1[2405]<=26'd1935091; ROM2[2405]<=26'd11272788; ROM3[2405]<=26'd9748624; ROM4[2405]<=26'd23452850;
ROM1[2406]<=26'd1938613; ROM2[2406]<=26'd11271551; ROM3[2406]<=26'd9742960; ROM4[2406]<=26'd23450626;
ROM1[2407]<=26'd1950665; ROM2[2407]<=26'd11272599; ROM3[2407]<=26'd9736866; ROM4[2407]<=26'd23449907;
ROM1[2408]<=26'd1955068; ROM2[2408]<=26'd11270664; ROM3[2408]<=26'd9729739; ROM4[2408]<=26'd23444968;
ROM1[2409]<=26'd1953136; ROM2[2409]<=26'd11273824; ROM3[2409]<=26'd9735791; ROM4[2409]<=26'd23448483;
ROM1[2410]<=26'd1947922; ROM2[2410]<=26'd11273727; ROM3[2410]<=26'd9742365; ROM4[2410]<=26'd23451904;
ROM1[2411]<=26'd1941257; ROM2[2411]<=26'd11271944; ROM3[2411]<=26'd9743819; ROM4[2411]<=26'd23451678;
ROM1[2412]<=26'd1936878; ROM2[2412]<=26'd11273082; ROM3[2412]<=26'd9744657; ROM4[2412]<=26'd23452370;
ROM1[2413]<=26'd1933522; ROM2[2413]<=26'd11272803; ROM3[2413]<=26'd9745245; ROM4[2413]<=26'd23452890;
ROM1[2414]<=26'd1936973; ROM2[2414]<=26'd11276022; ROM3[2414]<=26'd9744580; ROM4[2414]<=26'd23453960;
ROM1[2415]<=26'd1946617; ROM2[2415]<=26'd11278235; ROM3[2415]<=26'd9740231; ROM4[2415]<=26'd23454433;
ROM1[2416]<=26'd1959304; ROM2[2416]<=26'd11278756; ROM3[2416]<=26'd9736860; ROM4[2416]<=26'd23454510;
ROM1[2417]<=26'd1966070; ROM2[2417]<=26'd11283068; ROM3[2417]<=26'd9740879; ROM4[2417]<=26'd23459439;
ROM1[2418]<=26'd1960589; ROM2[2418]<=26'd11283613; ROM3[2418]<=26'd9744867; ROM4[2418]<=26'd23460656;
ROM1[2419]<=26'd1948943; ROM2[2419]<=26'd11277393; ROM3[2419]<=26'd9745061; ROM4[2419]<=26'd23456001;
ROM1[2420]<=26'd1942759; ROM2[2420]<=26'd11274948; ROM3[2420]<=26'd9745335; ROM4[2420]<=26'd23454987;
ROM1[2421]<=26'd1930804; ROM2[2421]<=26'd11269030; ROM3[2421]<=26'd9741147; ROM4[2421]<=26'd23449931;
ROM1[2422]<=26'd1932588; ROM2[2422]<=26'd11269378; ROM3[2422]<=26'd9742501; ROM4[2422]<=26'd23449875;
ROM1[2423]<=26'd1947796; ROM2[2423]<=26'd11276110; ROM3[2423]<=26'd9744505; ROM4[2423]<=26'd23454760;
ROM1[2424]<=26'd1959266; ROM2[2424]<=26'd11276526; ROM3[2424]<=26'd9741900; ROM4[2424]<=26'd23455320;
ROM1[2425]<=26'd1964453; ROM2[2425]<=26'd11278501; ROM3[2425]<=26'd9742819; ROM4[2425]<=26'd23458672;
ROM1[2426]<=26'd1964190; ROM2[2426]<=26'd11283938; ROM3[2426]<=26'd9749448; ROM4[2426]<=26'd23465728;
ROM1[2427]<=26'd1959441; ROM2[2427]<=26'd11285316; ROM3[2427]<=26'd9756103; ROM4[2427]<=26'd23467767;
ROM1[2428]<=26'd1950114; ROM2[2428]<=26'd11280740; ROM3[2428]<=26'd9752840; ROM4[2428]<=26'd23462408;
ROM1[2429]<=26'd1944535; ROM2[2429]<=26'd11279794; ROM3[2429]<=26'd9754880; ROM4[2429]<=26'd23462561;
ROM1[2430]<=26'd1943125; ROM2[2430]<=26'd11280772; ROM3[2430]<=26'd9756688; ROM4[2430]<=26'd23464035;
ROM1[2431]<=26'd1943382; ROM2[2431]<=26'd11277457; ROM3[2431]<=26'd9746691; ROM4[2431]<=26'd23458653;
ROM1[2432]<=26'd1958954; ROM2[2432]<=26'd11282258; ROM3[2432]<=26'd9743041; ROM4[2432]<=26'd23461672;
ROM1[2433]<=26'd1970830; ROM2[2433]<=26'd11286600; ROM3[2433]<=26'd9742173; ROM4[2433]<=26'd23464779;
ROM1[2434]<=26'd1963321; ROM2[2434]<=26'd11282469; ROM3[2434]<=26'd9737937; ROM4[2434]<=26'd23458635;
ROM1[2435]<=26'd1952973; ROM2[2435]<=26'd11277235; ROM3[2435]<=26'd9737749; ROM4[2435]<=26'd23454893;
ROM1[2436]<=26'd1948382; ROM2[2436]<=26'd11277017; ROM3[2436]<=26'd9742520; ROM4[2436]<=26'd23456594;
ROM1[2437]<=26'd1942498; ROM2[2437]<=26'd11277676; ROM3[2437]<=26'd9743782; ROM4[2437]<=26'd23456345;
ROM1[2438]<=26'd1938093; ROM2[2438]<=26'd11275648; ROM3[2438]<=26'd9744191; ROM4[2438]<=26'd23455549;
ROM1[2439]<=26'd1945012; ROM2[2439]<=26'd11280037; ROM3[2439]<=26'd9748585; ROM4[2439]<=26'd23459471;
ROM1[2440]<=26'd1954384; ROM2[2440]<=26'd11280759; ROM3[2440]<=26'd9745132; ROM4[2440]<=26'd23459994;
ROM1[2441]<=26'd1963033; ROM2[2441]<=26'd11279435; ROM3[2441]<=26'd9738644; ROM4[2441]<=26'd23456825;
ROM1[2442]<=26'd1961659; ROM2[2442]<=26'd11280094; ROM3[2442]<=26'd9738681; ROM4[2442]<=26'd23456271;
ROM1[2443]<=26'd1954707; ROM2[2443]<=26'd11279880; ROM3[2443]<=26'd9741994; ROM4[2443]<=26'd23458601;
ROM1[2444]<=26'd1946025; ROM2[2444]<=26'd11278775; ROM3[2444]<=26'd9744475; ROM4[2444]<=26'd23458037;
ROM1[2445]<=26'd1937199; ROM2[2445]<=26'd11275325; ROM3[2445]<=26'd9742422; ROM4[2445]<=26'd23454763;
ROM1[2446]<=26'd1931570; ROM2[2446]<=26'd11272946; ROM3[2446]<=26'd9740968; ROM4[2446]<=26'd23453045;
ROM1[2447]<=26'd1932376; ROM2[2447]<=26'd11273268; ROM3[2447]<=26'd9740465; ROM4[2447]<=26'd23452620;
ROM1[2448]<=26'd1940425; ROM2[2448]<=26'd11274861; ROM3[2448]<=26'd9736449; ROM4[2448]<=26'd23452353;
ROM1[2449]<=26'd1955104; ROM2[2449]<=26'd11279107; ROM3[2449]<=26'd9731854; ROM4[2449]<=26'd23454861;
ROM1[2450]<=26'd1957589; ROM2[2450]<=26'd11280179; ROM3[2450]<=26'd9730549; ROM4[2450]<=26'd23454606;
ROM1[2451]<=26'd1951739; ROM2[2451]<=26'd11278994; ROM3[2451]<=26'd9733137; ROM4[2451]<=26'd23454443;
ROM1[2452]<=26'd1947787; ROM2[2452]<=26'd11278942; ROM3[2452]<=26'd9737526; ROM4[2452]<=26'd23456766;
ROM1[2453]<=26'd1941699; ROM2[2453]<=26'd11275810; ROM3[2453]<=26'd9738498; ROM4[2453]<=26'd23455150;
ROM1[2454]<=26'd1936409; ROM2[2454]<=26'd11276895; ROM3[2454]<=26'd9741725; ROM4[2454]<=26'd23456776;
ROM1[2455]<=26'd1936207; ROM2[2455]<=26'd11281557; ROM3[2455]<=26'd9744348; ROM4[2455]<=26'd23459499;
ROM1[2456]<=26'd1939932; ROM2[2456]<=26'd11281972; ROM3[2456]<=26'd9741878; ROM4[2456]<=26'd23457405;
ROM1[2457]<=26'd1949357; ROM2[2457]<=26'd11280660; ROM3[2457]<=26'd9735300; ROM4[2457]<=26'd23453859;
ROM1[2458]<=26'd1958888; ROM2[2458]<=26'd11280527; ROM3[2458]<=26'd9732348; ROM4[2458]<=26'd23454537;
ROM1[2459]<=26'd1956518; ROM2[2459]<=26'd11281794; ROM3[2459]<=26'd9734006; ROM4[2459]<=26'd23455279;
ROM1[2460]<=26'd1952180; ROM2[2460]<=26'd11285219; ROM3[2460]<=26'd9739611; ROM4[2460]<=26'd23458061;
ROM1[2461]<=26'd1952881; ROM2[2461]<=26'd11289859; ROM3[2461]<=26'd9747838; ROM4[2461]<=26'd23463557;
ROM1[2462]<=26'd1946310; ROM2[2462]<=26'd11286358; ROM3[2462]<=26'd9747136; ROM4[2462]<=26'd23459771;
ROM1[2463]<=26'd1940959; ROM2[2463]<=26'd11282002; ROM3[2463]<=26'd9746970; ROM4[2463]<=26'd23458799;
ROM1[2464]<=26'd1940506; ROM2[2464]<=26'd11278919; ROM3[2464]<=26'd9743663; ROM4[2464]<=26'd23456625;
ROM1[2465]<=26'd1944184; ROM2[2465]<=26'd11274664; ROM3[2465]<=26'd9736318; ROM4[2465]<=26'd23450461;
ROM1[2466]<=26'd1955610; ROM2[2466]<=26'd11277220; ROM3[2466]<=26'd9734256; ROM4[2466]<=26'd23451220;
ROM1[2467]<=26'd1955224; ROM2[2467]<=26'd11278631; ROM3[2467]<=26'd9733612; ROM4[2467]<=26'd23451564;
ROM1[2468]<=26'd1949454; ROM2[2468]<=26'd11277782; ROM3[2468]<=26'd9736313; ROM4[2468]<=26'd23452088;
ROM1[2469]<=26'd1945731; ROM2[2469]<=26'd11278444; ROM3[2469]<=26'd9743536; ROM4[2469]<=26'd23455640;
ROM1[2470]<=26'd1942869; ROM2[2470]<=26'd11279377; ROM3[2470]<=26'd9745551; ROM4[2470]<=26'd23456983;
ROM1[2471]<=26'd1936777; ROM2[2471]<=26'd11277825; ROM3[2471]<=26'd9746563; ROM4[2471]<=26'd23454357;
ROM1[2472]<=26'd1937802; ROM2[2472]<=26'd11278711; ROM3[2472]<=26'd9747710; ROM4[2472]<=26'd23455714;
ROM1[2473]<=26'd1946638; ROM2[2473]<=26'd11280201; ROM3[2473]<=26'd9742810; ROM4[2473]<=26'd23456174;
ROM1[2474]<=26'd1956016; ROM2[2474]<=26'd11278012; ROM3[2474]<=26'd9734782; ROM4[2474]<=26'd23451624;
ROM1[2475]<=26'd1961039; ROM2[2475]<=26'd11278796; ROM3[2475]<=26'd9733693; ROM4[2475]<=26'd23453461;
ROM1[2476]<=26'd1958374; ROM2[2476]<=26'd11281003; ROM3[2476]<=26'd9738925; ROM4[2476]<=26'd23455351;
ROM1[2477]<=26'd1952075; ROM2[2477]<=26'd11280935; ROM3[2477]<=26'd9744347; ROM4[2477]<=26'd23455727;
ROM1[2478]<=26'd1945428; ROM2[2478]<=26'd11277330; ROM3[2478]<=26'd9744972; ROM4[2478]<=26'd23455178;
ROM1[2479]<=26'd1931039; ROM2[2479]<=26'd11267103; ROM3[2479]<=26'd9738604; ROM4[2479]<=26'd23446923;
ROM1[2480]<=26'd1925278; ROM2[2480]<=26'd11263396; ROM3[2480]<=26'd9735726; ROM4[2480]<=26'd23443248;
ROM1[2481]<=26'd1931417; ROM2[2481]<=26'd11266325; ROM3[2481]<=26'd9731908; ROM4[2481]<=26'd23443051;
ROM1[2482]<=26'd1947549; ROM2[2482]<=26'd11271015; ROM3[2482]<=26'd9729591; ROM4[2482]<=26'd23445667;
ROM1[2483]<=26'd1959456; ROM2[2483]<=26'd11273905; ROM3[2483]<=26'd9728665; ROM4[2483]<=26'd23447994;
ROM1[2484]<=26'd1953493; ROM2[2484]<=26'd11272527; ROM3[2484]<=26'd9725805; ROM4[2484]<=26'd23445291;
ROM1[2485]<=26'd1944617; ROM2[2485]<=26'd11270689; ROM3[2485]<=26'd9728256; ROM4[2485]<=26'd23442415;
ROM1[2486]<=26'd1940261; ROM2[2486]<=26'd11272428; ROM3[2486]<=26'd9734490; ROM4[2486]<=26'd23445054;
ROM1[2487]<=26'd1940082; ROM2[2487]<=26'd11277234; ROM3[2487]<=26'd9740417; ROM4[2487]<=26'd23449276;
ROM1[2488]<=26'd1940768; ROM2[2488]<=26'd11280989; ROM3[2488]<=26'd9747406; ROM4[2488]<=26'd23453186;
ROM1[2489]<=26'd1943640; ROM2[2489]<=26'd11281283; ROM3[2489]<=26'd9748841; ROM4[2489]<=26'd23455187;
ROM1[2490]<=26'd1946824; ROM2[2490]<=26'd11275131; ROM3[2490]<=26'd9737499; ROM4[2490]<=26'd23446820;
ROM1[2491]<=26'd1951912; ROM2[2491]<=26'd11269513; ROM3[2491]<=26'd9727527; ROM4[2491]<=26'd23439942;
ROM1[2492]<=26'd1950294; ROM2[2492]<=26'd11266884; ROM3[2492]<=26'd9726680; ROM4[2492]<=26'd23438461;
ROM1[2493]<=26'd1943267; ROM2[2493]<=26'd11267009; ROM3[2493]<=26'd9727865; ROM4[2493]<=26'd23439709;
ROM1[2494]<=26'd1946036; ROM2[2494]<=26'd11276888; ROM3[2494]<=26'd9739461; ROM4[2494]<=26'd23450411;
ROM1[2495]<=26'd1950416; ROM2[2495]<=26'd11284374; ROM3[2495]<=26'd9748852; ROM4[2495]<=26'd23458791;
ROM1[2496]<=26'd1940832; ROM2[2496]<=26'd11279998; ROM3[2496]<=26'd9745670; ROM4[2496]<=26'd23455044;
ROM1[2497]<=26'd1930400; ROM2[2497]<=26'd11269249; ROM3[2497]<=26'd9734364; ROM4[2497]<=26'd23443392;
ROM1[2498]<=26'd1934002; ROM2[2498]<=26'd11263223; ROM3[2498]<=26'd9727034; ROM4[2498]<=26'd23438420;
ROM1[2499]<=26'd1948038; ROM2[2499]<=26'd11269117; ROM3[2499]<=26'd9723860; ROM4[2499]<=26'd23440952;
ROM1[2500]<=26'd1956529; ROM2[2500]<=26'd11274315; ROM3[2500]<=26'd9722805; ROM4[2500]<=26'd23443822;
ROM1[2501]<=26'd1951607; ROM2[2501]<=26'd11272258; ROM3[2501]<=26'd9725640; ROM4[2501]<=26'd23445072;
ROM1[2502]<=26'd1942279; ROM2[2502]<=26'd11271362; ROM3[2502]<=26'd9729109; ROM4[2502]<=26'd23444790;
ROM1[2503]<=26'd1937573; ROM2[2503]<=26'd11271599; ROM3[2503]<=26'd9732569; ROM4[2503]<=26'd23446862;
ROM1[2504]<=26'd1927743; ROM2[2504]<=26'd11268964; ROM3[2504]<=26'd9733072; ROM4[2504]<=26'd23446621;
ROM1[2505]<=26'd1928900; ROM2[2505]<=26'd11271640; ROM3[2505]<=26'd9737303; ROM4[2505]<=26'd23447646;
ROM1[2506]<=26'd1937063; ROM2[2506]<=26'd11274436; ROM3[2506]<=26'd9736945; ROM4[2506]<=26'd23449429;
ROM1[2507]<=26'd1952750; ROM2[2507]<=26'd11278189; ROM3[2507]<=26'd9735759; ROM4[2507]<=26'd23453055;
ROM1[2508]<=26'd1963258; ROM2[2508]<=26'd11279497; ROM3[2508]<=26'd9733616; ROM4[2508]<=26'd23454070;
ROM1[2509]<=26'd1953169; ROM2[2509]<=26'd11274468; ROM3[2509]<=26'd9727028; ROM4[2509]<=26'd23448846;
ROM1[2510]<=26'd1944835; ROM2[2510]<=26'd11273223; ROM3[2510]<=26'd9730322; ROM4[2510]<=26'd23447535;
ROM1[2511]<=26'd1939203; ROM2[2511]<=26'd11272072; ROM3[2511]<=26'd9734741; ROM4[2511]<=26'd23448453;
ROM1[2512]<=26'd1933174; ROM2[2512]<=26'd11269991; ROM3[2512]<=26'd9737864; ROM4[2512]<=26'd23448358;
ROM1[2513]<=26'd1934937; ROM2[2513]<=26'd11273011; ROM3[2513]<=26'd9745237; ROM4[2513]<=26'd23453192;
ROM1[2514]<=26'd1941351; ROM2[2514]<=26'd11276680; ROM3[2514]<=26'd9747397; ROM4[2514]<=26'd23457498;
ROM1[2515]<=26'd1949868; ROM2[2515]<=26'd11277666; ROM3[2515]<=26'd9743171; ROM4[2515]<=26'd23455999;
ROM1[2516]<=26'd1963877; ROM2[2516]<=26'd11280763; ROM3[2516]<=26'd9739769; ROM4[2516]<=26'd23458053;
ROM1[2517]<=26'd1969394; ROM2[2517]<=26'd11285970; ROM3[2517]<=26'd9743861; ROM4[2517]<=26'd23463587;
ROM1[2518]<=26'd1960669; ROM2[2518]<=26'd11283363; ROM3[2518]<=26'd9744233; ROM4[2518]<=26'd23462113;
ROM1[2519]<=26'd1947304; ROM2[2519]<=26'd11275111; ROM3[2519]<=26'd9739918; ROM4[2519]<=26'd23456046;
ROM1[2520]<=26'd1942733; ROM2[2520]<=26'd11273946; ROM3[2520]<=26'd9741856; ROM4[2520]<=26'd23455294;
ROM1[2521]<=26'd1938131; ROM2[2521]<=26'd11274876; ROM3[2521]<=26'd9746656; ROM4[2521]<=26'd23457955;
ROM1[2522]<=26'd1937309; ROM2[2522]<=26'd11275943; ROM3[2522]<=26'd9747774; ROM4[2522]<=26'd23458992;
ROM1[2523]<=26'd1946928; ROM2[2523]<=26'd11279569; ROM3[2523]<=26'd9745586; ROM4[2523]<=26'd23458152;
ROM1[2524]<=26'd1959602; ROM2[2524]<=26'd11279354; ROM3[2524]<=26'd9741444; ROM4[2524]<=26'd23457698;
ROM1[2525]<=26'd1963318; ROM2[2525]<=26'd11279153; ROM3[2525]<=26'd9739237; ROM4[2525]<=26'd23458121;
ROM1[2526]<=26'd1957474; ROM2[2526]<=26'd11278787; ROM3[2526]<=26'd9743051; ROM4[2526]<=26'd23460309;
ROM1[2527]<=26'd1957040; ROM2[2527]<=26'd11283222; ROM3[2527]<=26'd9754672; ROM4[2527]<=26'd23468629;
ROM1[2528]<=26'd1960274; ROM2[2528]<=26'd11289312; ROM3[2528]<=26'd9764993; ROM4[2528]<=26'd23475211;
ROM1[2529]<=26'd1951795; ROM2[2529]<=26'd11284478; ROM3[2529]<=26'd9765001; ROM4[2529]<=26'd23471601;
ROM1[2530]<=26'd1948603; ROM2[2530]<=26'd11283023; ROM3[2530]<=26'd9763072; ROM4[2530]<=26'd23469208;
ROM1[2531]<=26'd1949783; ROM2[2531]<=26'd11279410; ROM3[2531]<=26'd9756791; ROM4[2531]<=26'd23464651;
ROM1[2532]<=26'd1958855; ROM2[2532]<=26'd11278872; ROM3[2532]<=26'd9750396; ROM4[2532]<=26'd23464378;
ROM1[2533]<=26'd1974291; ROM2[2533]<=26'd11286320; ROM3[2533]<=26'd9751472; ROM4[2533]<=26'd23470507;
ROM1[2534]<=26'd1976334; ROM2[2534]<=26'd11288172; ROM3[2534]<=26'd9752185; ROM4[2534]<=26'd23472034;
ROM1[2535]<=26'd1969347; ROM2[2535]<=26'd11287828; ROM3[2535]<=26'd9756347; ROM4[2535]<=26'd23473139;
ROM1[2536]<=26'd1962969; ROM2[2536]<=26'd11287151; ROM3[2536]<=26'd9758654; ROM4[2536]<=26'd23471933;
ROM1[2537]<=26'd1957105; ROM2[2537]<=26'd11287020; ROM3[2537]<=26'd9758484; ROM4[2537]<=26'd23470357;
ROM1[2538]<=26'd1955184; ROM2[2538]<=26'd11287717; ROM3[2538]<=26'd9761864; ROM4[2538]<=26'd23472125;
ROM1[2539]<=26'd1959579; ROM2[2539]<=26'd11288117; ROM3[2539]<=26'd9758542; ROM4[2539]<=26'd23471347;
ROM1[2540]<=26'd1965619; ROM2[2540]<=26'd11286117; ROM3[2540]<=26'd9748500; ROM4[2540]<=26'd23465925;
ROM1[2541]<=26'd1977434; ROM2[2541]<=26'd11288515; ROM3[2541]<=26'd9745249; ROM4[2541]<=26'd23467210;
ROM1[2542]<=26'd1981094; ROM2[2542]<=26'd11292293; ROM3[2542]<=26'd9746327; ROM4[2542]<=26'd23469677;
ROM1[2543]<=26'd1974288; ROM2[2543]<=26'd11291844; ROM3[2543]<=26'd9748633; ROM4[2543]<=26'd23469131;
ROM1[2544]<=26'd1975717; ROM2[2544]<=26'd11301300; ROM3[2544]<=26'd9762027; ROM4[2544]<=26'd23479145;
ROM1[2545]<=26'd1972331; ROM2[2545]<=26'd11303208; ROM3[2545]<=26'd9766533; ROM4[2545]<=26'd23481337;
ROM1[2546]<=26'd1958070; ROM2[2546]<=26'd11293419; ROM3[2546]<=26'd9761011; ROM4[2546]<=26'd23473240;
ROM1[2547]<=26'd1955558; ROM2[2547]<=26'd11290443; ROM3[2547]<=26'd9759085; ROM4[2547]<=26'd23470587;
ROM1[2548]<=26'd1955632; ROM2[2548]<=26'd11282343; ROM3[2548]<=26'd9747162; ROM4[2548]<=26'd23461873;
ROM1[2549]<=26'd1968205; ROM2[2549]<=26'd11283214; ROM3[2549]<=26'd9740275; ROM4[2549]<=26'd23462176;
ROM1[2550]<=26'd1974503; ROM2[2550]<=26'd11285185; ROM3[2550]<=26'd9740724; ROM4[2550]<=26'd23463896;
ROM1[2551]<=26'd1970304; ROM2[2551]<=26'd11285023; ROM3[2551]<=26'd9743201; ROM4[2551]<=26'd23464542;
ROM1[2552]<=26'd1966233; ROM2[2552]<=26'd11286916; ROM3[2552]<=26'd9749162; ROM4[2552]<=26'd23468136;
ROM1[2553]<=26'd1961001; ROM2[2553]<=26'd11286394; ROM3[2553]<=26'd9753403; ROM4[2553]<=26'd23468791;
ROM1[2554]<=26'd1956358; ROM2[2554]<=26'd11288107; ROM3[2554]<=26'd9758484; ROM4[2554]<=26'd23469595;
ROM1[2555]<=26'd1952120; ROM2[2555]<=26'd11285764; ROM3[2555]<=26'd9755718; ROM4[2555]<=26'd23466702;
ROM1[2556]<=26'd1957011; ROM2[2556]<=26'd11285747; ROM3[2556]<=26'd9750712; ROM4[2556]<=26'd23464500;
ROM1[2557]<=26'd1969618; ROM2[2557]<=26'd11287121; ROM3[2557]<=26'd9744221; ROM4[2557]<=26'd23463082;
ROM1[2558]<=26'd1975905; ROM2[2558]<=26'd11285964; ROM3[2558]<=26'd9739057; ROM4[2558]<=26'd23462704;
ROM1[2559]<=26'd1974092; ROM2[2559]<=26'd11287917; ROM3[2559]<=26'd9740390; ROM4[2559]<=26'd23464406;
ROM1[2560]<=26'd1971682; ROM2[2560]<=26'd11293176; ROM3[2560]<=26'd9746374; ROM4[2560]<=26'd23467787;
ROM1[2561]<=26'd1970871; ROM2[2561]<=26'd11297994; ROM3[2561]<=26'd9756415; ROM4[2561]<=26'd23472694;
ROM1[2562]<=26'd1960082; ROM2[2562]<=26'd11293701; ROM3[2562]<=26'd9755382; ROM4[2562]<=26'd23470209;
ROM1[2563]<=26'd1951312; ROM2[2563]<=26'd11288925; ROM3[2563]<=26'd9753543; ROM4[2563]<=26'd23465960;
ROM1[2564]<=26'd1950743; ROM2[2564]<=26'd11284804; ROM3[2564]<=26'd9752480; ROM4[2564]<=26'd23463318;
ROM1[2565]<=26'd1956000; ROM2[2565]<=26'd11281798; ROM3[2565]<=26'd9744214; ROM4[2565]<=26'd23460067;
ROM1[2566]<=26'd1969766; ROM2[2566]<=26'd11287607; ROM3[2566]<=26'd9740065; ROM4[2566]<=26'd23462554;
ROM1[2567]<=26'd1973561; ROM2[2567]<=26'd11291055; ROM3[2567]<=26'd9743917; ROM4[2567]<=26'd23466661;
ROM1[2568]<=26'd1967851; ROM2[2568]<=26'd11290166; ROM3[2568]<=26'd9747540; ROM4[2568]<=26'd23467364;
ROM1[2569]<=26'd1962839; ROM2[2569]<=26'd11289830; ROM3[2569]<=26'd9751938; ROM4[2569]<=26'd23467450;
ROM1[2570]<=26'd1959838; ROM2[2570]<=26'd11291419; ROM3[2570]<=26'd9757541; ROM4[2570]<=26'd23469608;
ROM1[2571]<=26'd1953821; ROM2[2571]<=26'd11291075; ROM3[2571]<=26'd9762418; ROM4[2571]<=26'd23469728;
ROM1[2572]<=26'd1948799; ROM2[2572]<=26'd11285883; ROM3[2572]<=26'd9758592; ROM4[2572]<=26'd23465010;
ROM1[2573]<=26'd1953742; ROM2[2573]<=26'd11285031; ROM3[2573]<=26'd9752021; ROM4[2573]<=26'd23463752;
ROM1[2574]<=26'd1970100; ROM2[2574]<=26'd11287550; ROM3[2574]<=26'd9750396; ROM4[2574]<=26'd23465103;
ROM1[2575]<=26'd1977085; ROM2[2575]<=26'd11290586; ROM3[2575]<=26'd9750051; ROM4[2575]<=26'd23467597;
ROM1[2576]<=26'd1974862; ROM2[2576]<=26'd11293114; ROM3[2576]<=26'd9753270; ROM4[2576]<=26'd23470997;
ROM1[2577]<=26'd1966207; ROM2[2577]<=26'd11291070; ROM3[2577]<=26'd9755361; ROM4[2577]<=26'd23468858;
ROM1[2578]<=26'd1958955; ROM2[2578]<=26'd11290137; ROM3[2578]<=26'd9755540; ROM4[2578]<=26'd23468042;
ROM1[2579]<=26'd1949934; ROM2[2579]<=26'd11287082; ROM3[2579]<=26'd9754388; ROM4[2579]<=26'd23466387;
ROM1[2580]<=26'd1945022; ROM2[2580]<=26'd11284671; ROM3[2580]<=26'd9751862; ROM4[2580]<=26'd23463979;
ROM1[2581]<=26'd1953345; ROM2[2581]<=26'd11286878; ROM3[2581]<=26'd9751011; ROM4[2581]<=26'd23465597;
ROM1[2582]<=26'd1971959; ROM2[2582]<=26'd11291623; ROM3[2582]<=26'd9750675; ROM4[2582]<=26'd23468777;
ROM1[2583]<=26'd1984032; ROM2[2583]<=26'd11294441; ROM3[2583]<=26'd9748549; ROM4[2583]<=26'd23472059;
ROM1[2584]<=26'd1981070; ROM2[2584]<=26'd11296028; ROM3[2584]<=26'd9751302; ROM4[2584]<=26'd23474267;
ROM1[2585]<=26'd1974990; ROM2[2585]<=26'd11296865; ROM3[2585]<=26'd9756149; ROM4[2585]<=26'd23476392;
ROM1[2586]<=26'd1970328; ROM2[2586]<=26'd11297168; ROM3[2586]<=26'd9761503; ROM4[2586]<=26'd23479720;
ROM1[2587]<=26'd1964902; ROM2[2587]<=26'd11296177; ROM3[2587]<=26'd9765252; ROM4[2587]<=26'd23479294;
ROM1[2588]<=26'd1958922; ROM2[2588]<=26'd11295322; ROM3[2588]<=26'd9766516; ROM4[2588]<=26'd23478541;
ROM1[2589]<=26'd1958084; ROM2[2589]<=26'd11292860; ROM3[2589]<=26'd9762656; ROM4[2589]<=26'd23476123;
ROM1[2590]<=26'd1965052; ROM2[2590]<=26'd11289597; ROM3[2590]<=26'd9753658; ROM4[2590]<=26'd23470753;
ROM1[2591]<=26'd1975480; ROM2[2591]<=26'd11291424; ROM3[2591]<=26'd9747505; ROM4[2591]<=26'd23469344;
ROM1[2592]<=26'd1974880; ROM2[2592]<=26'd11290547; ROM3[2592]<=26'd9744507; ROM4[2592]<=26'd23467438;
ROM1[2593]<=26'd1967227; ROM2[2593]<=26'd11288951; ROM3[2593]<=26'd9745537; ROM4[2593]<=26'd23466952;
ROM1[2594]<=26'd1959005; ROM2[2594]<=26'd11288869; ROM3[2594]<=26'd9746946; ROM4[2594]<=26'd23466956;
ROM1[2595]<=26'd1958479; ROM2[2595]<=26'd11294388; ROM3[2595]<=26'd9752836; ROM4[2595]<=26'd23471193;
ROM1[2596]<=26'd1956254; ROM2[2596]<=26'd11297559; ROM3[2596]<=26'd9755852; ROM4[2596]<=26'd23473278;
ROM1[2597]<=26'd1953442; ROM2[2597]<=26'd11295370; ROM3[2597]<=26'd9750213; ROM4[2597]<=26'd23467733;
ROM1[2598]<=26'd1960006; ROM2[2598]<=26'd11294360; ROM3[2598]<=26'd9745469; ROM4[2598]<=26'd23464722;
ROM1[2599]<=26'd1967382; ROM2[2599]<=26'd11290297; ROM3[2599]<=26'd9735501; ROM4[2599]<=26'd23459352;
ROM1[2600]<=26'd1966626; ROM2[2600]<=26'd11285950; ROM3[2600]<=26'd9731233; ROM4[2600]<=26'd23456385;
ROM1[2601]<=26'd1964029; ROM2[2601]<=26'd11286513; ROM3[2601]<=26'd9737894; ROM4[2601]<=26'd23459205;
ROM1[2602]<=26'd1958592; ROM2[2602]<=26'd11288710; ROM3[2602]<=26'd9745499; ROM4[2602]<=26'd23460958;
ROM1[2603]<=26'd1951594; ROM2[2603]<=26'd11285282; ROM3[2603]<=26'd9746036; ROM4[2603]<=26'd23459622;
ROM1[2604]<=26'd1949179; ROM2[2604]<=26'd11287335; ROM3[2604]<=26'd9750431; ROM4[2604]<=26'd23462439;
ROM1[2605]<=26'd1951612; ROM2[2605]<=26'd11290237; ROM3[2605]<=26'd9757506; ROM4[2605]<=26'd23466704;
ROM1[2606]<=26'd1955667; ROM2[2606]<=26'd11290712; ROM3[2606]<=26'd9755714; ROM4[2606]<=26'd23467605;
ROM1[2607]<=26'd1965826; ROM2[2607]<=26'd11290633; ROM3[2607]<=26'd9750434; ROM4[2607]<=26'd23467767;
ROM1[2608]<=26'd1975350; ROM2[2608]<=26'd11292670; ROM3[2608]<=26'd9748343; ROM4[2608]<=26'd23468789;
ROM1[2609]<=26'd1976316; ROM2[2609]<=26'd11299715; ROM3[2609]<=26'd9754046; ROM4[2609]<=26'd23475210;
ROM1[2610]<=26'd1968345; ROM2[2610]<=26'd11296751; ROM3[2610]<=26'd9756962; ROM4[2610]<=26'd23475885;
ROM1[2611]<=26'd1954285; ROM2[2611]<=26'd11287430; ROM3[2611]<=26'd9752983; ROM4[2611]<=26'd23468342;
ROM1[2612]<=26'd1945317; ROM2[2612]<=26'd11285055; ROM3[2612]<=26'd9754033; ROM4[2612]<=26'd23467043;
ROM1[2613]<=26'd1938210; ROM2[2613]<=26'd11280083; ROM3[2613]<=26'd9750536; ROM4[2613]<=26'd23462194;
ROM1[2614]<=26'd1943147; ROM2[2614]<=26'd11282889; ROM3[2614]<=26'd9749587; ROM4[2614]<=26'd23461213;
ROM1[2615]<=26'd1961764; ROM2[2615]<=26'd11294980; ROM3[2615]<=26'd9755705; ROM4[2615]<=26'd23468840;
ROM1[2616]<=26'd1967389; ROM2[2616]<=26'd11289177; ROM3[2616]<=26'd9745314; ROM4[2616]<=26'd23462117;
ROM1[2617]<=26'd1962632; ROM2[2617]<=26'd11282575; ROM3[2617]<=26'd9737039; ROM4[2617]<=26'd23455026;
ROM1[2618]<=26'd1957714; ROM2[2618]<=26'd11281092; ROM3[2618]<=26'd9737854; ROM4[2618]<=26'd23453701;
ROM1[2619]<=26'd1952335; ROM2[2619]<=26'd11280630; ROM3[2619]<=26'd9739996; ROM4[2619]<=26'd23452986;
ROM1[2620]<=26'd1951706; ROM2[2620]<=26'd11285161; ROM3[2620]<=26'd9745599; ROM4[2620]<=26'd23456877;
ROM1[2621]<=26'd1944633; ROM2[2621]<=26'd11284274; ROM3[2621]<=26'd9748364; ROM4[2621]<=26'd23456928;
ROM1[2622]<=26'd1943165; ROM2[2622]<=26'd11283599; ROM3[2622]<=26'd9748967; ROM4[2622]<=26'd23458014;
ROM1[2623]<=26'd1954131; ROM2[2623]<=26'd11285821; ROM3[2623]<=26'd9746529; ROM4[2623]<=26'd23460120;
ROM1[2624]<=26'd1968815; ROM2[2624]<=26'd11285775; ROM3[2624]<=26'd9741982; ROM4[2624]<=26'd23459403;
ROM1[2625]<=26'd1973310; ROM2[2625]<=26'd11286302; ROM3[2625]<=26'd9739965; ROM4[2625]<=26'd23459232;
ROM1[2626]<=26'd1965911; ROM2[2626]<=26'd11284642; ROM3[2626]<=26'd9740955; ROM4[2626]<=26'd23457624;
ROM1[2627]<=26'd1959266; ROM2[2627]<=26'd11282633; ROM3[2627]<=26'd9745454; ROM4[2627]<=26'd23457681;
ROM1[2628]<=26'd1959018; ROM2[2628]<=26'd11287877; ROM3[2628]<=26'd9752648; ROM4[2628]<=26'd23464157;
ROM1[2629]<=26'd1952316; ROM2[2629]<=26'd11286834; ROM3[2629]<=26'd9754506; ROM4[2629]<=26'd23463120;
ROM1[2630]<=26'd1945135; ROM2[2630]<=26'd11282419; ROM3[2630]<=26'd9747352; ROM4[2630]<=26'd23456530;
ROM1[2631]<=26'd1950255; ROM2[2631]<=26'd11283595; ROM3[2631]<=26'd9743339; ROM4[2631]<=26'd23455833;
ROM1[2632]<=26'd1961223; ROM2[2632]<=26'd11283320; ROM3[2632]<=26'd9738020; ROM4[2632]<=26'd23454216;
ROM1[2633]<=26'd1967798; ROM2[2633]<=26'd11284074; ROM3[2633]<=26'd9733745; ROM4[2633]<=26'd23453573;
ROM1[2634]<=26'd1962436; ROM2[2634]<=26'd11283320; ROM3[2634]<=26'd9734192; ROM4[2634]<=26'd23453169;
ROM1[2635]<=26'd1948918; ROM2[2635]<=26'd11278490; ROM3[2635]<=26'd9732952; ROM4[2635]<=26'd23447901;
ROM1[2636]<=26'd1943854; ROM2[2636]<=26'd11280713; ROM3[2636]<=26'd9737393; ROM4[2636]<=26'd23450286;
ROM1[2637]<=26'd1943555; ROM2[2637]<=26'd11283962; ROM3[2637]<=26'd9744706; ROM4[2637]<=26'd23456696;
ROM1[2638]<=26'd1941004; ROM2[2638]<=26'd11283371; ROM3[2638]<=26'd9747913; ROM4[2638]<=26'd23458705;
ROM1[2639]<=26'd1944428; ROM2[2639]<=26'd11284502; ROM3[2639]<=26'd9749186; ROM4[2639]<=26'd23461309;
ROM1[2640]<=26'd1952254; ROM2[2640]<=26'd11282873; ROM3[2640]<=26'd9743548; ROM4[2640]<=26'd23457419;
ROM1[2641]<=26'd1962613; ROM2[2641]<=26'd11282864; ROM3[2641]<=26'd9735838; ROM4[2641]<=26'd23454874;
ROM1[2642]<=26'd1966747; ROM2[2642]<=26'd11284420; ROM3[2642]<=26'd9735907; ROM4[2642]<=26'd23457587;
ROM1[2643]<=26'd1962140; ROM2[2643]<=26'd11285505; ROM3[2643]<=26'd9739204; ROM4[2643]<=26'd23459816;
ROM1[2644]<=26'd1956331; ROM2[2644]<=26'd11286425; ROM3[2644]<=26'd9742629; ROM4[2644]<=26'd23461188;
ROM1[2645]<=26'd1953779; ROM2[2645]<=26'd11287116; ROM3[2645]<=26'd9746649; ROM4[2645]<=26'd23463862;
ROM1[2646]<=26'd1948915; ROM2[2646]<=26'd11288258; ROM3[2646]<=26'd9747981; ROM4[2646]<=26'd23464346;
ROM1[2647]<=26'd1948534; ROM2[2647]<=26'd11288474; ROM3[2647]<=26'd9746028; ROM4[2647]<=26'd23462494;
ROM1[2648]<=26'd1957224; ROM2[2648]<=26'd11290354; ROM3[2648]<=26'd9743693; ROM4[2648]<=26'd23462144;
ROM1[2649]<=26'd1966273; ROM2[2649]<=26'd11290367; ROM3[2649]<=26'd9734835; ROM4[2649]<=26'd23459021;
ROM1[2650]<=26'd1964660; ROM2[2650]<=26'd11285853; ROM3[2650]<=26'd9730651; ROM4[2650]<=26'd23456162;
ROM1[2651]<=26'd1960513; ROM2[2651]<=26'd11285549; ROM3[2651]<=26'd9734588; ROM4[2651]<=26'd23459766;
ROM1[2652]<=26'd1953689; ROM2[2652]<=26'd11284901; ROM3[2652]<=26'd9737546; ROM4[2652]<=26'd23460475;
ROM1[2653]<=26'd1947640; ROM2[2653]<=26'd11284299; ROM3[2653]<=26'd9740970; ROM4[2653]<=26'd23461383;
ROM1[2654]<=26'd1942293; ROM2[2654]<=26'd11286570; ROM3[2654]<=26'd9745817; ROM4[2654]<=26'd23464584;
ROM1[2655]<=26'd1943305; ROM2[2655]<=26'd11289885; ROM3[2655]<=26'd9750338; ROM4[2655]<=26'd23465715;
ROM1[2656]<=26'd1951637; ROM2[2656]<=26'd11291872; ROM3[2656]<=26'd9749435; ROM4[2656]<=26'd23466842;
ROM1[2657]<=26'd1961014; ROM2[2657]<=26'd11291390; ROM3[2657]<=26'd9742120; ROM4[2657]<=26'd23464029;
ROM1[2658]<=26'd1973479; ROM2[2658]<=26'd11296864; ROM3[2658]<=26'd9742143; ROM4[2658]<=26'd23467552;
ROM1[2659]<=26'd1970989; ROM2[2659]<=26'd11296181; ROM3[2659]<=26'd9742760; ROM4[2659]<=26'd23467819;
ROM1[2660]<=26'd1954507; ROM2[2660]<=26'd11284550; ROM3[2660]<=26'd9737034; ROM4[2660]<=26'd23458848;
ROM1[2661]<=26'd1948508; ROM2[2661]<=26'd11283509; ROM3[2661]<=26'd9740915; ROM4[2661]<=26'd23459022;
ROM1[2662]<=26'd1944326; ROM2[2662]<=26'd11284152; ROM3[2662]<=26'd9743663; ROM4[2662]<=26'd23458888;
ROM1[2663]<=26'd1938920; ROM2[2663]<=26'd11282739; ROM3[2663]<=26'd9743031; ROM4[2663]<=26'd23456416;
ROM1[2664]<=26'd1944954; ROM2[2664]<=26'd11287559; ROM3[2664]<=26'd9746054; ROM4[2664]<=26'd23460132;
ROM1[2665]<=26'd1960156; ROM2[2665]<=26'd11292026; ROM3[2665]<=26'd9745298; ROM4[2665]<=26'd23462789;
ROM1[2666]<=26'd1972545; ROM2[2666]<=26'd11293206; ROM3[2666]<=26'd9741245; ROM4[2666]<=26'd23463173;
ROM1[2667]<=26'd1973629; ROM2[2667]<=26'd11293987; ROM3[2667]<=26'd9742936; ROM4[2667]<=26'd23466163;
ROM1[2668]<=26'd1968989; ROM2[2668]<=26'd11295687; ROM3[2668]<=26'd9749061; ROM4[2668]<=26'd23469625;
ROM1[2669]<=26'd1958727; ROM2[2669]<=26'd11290968; ROM3[2669]<=26'd9751217; ROM4[2669]<=26'd23466179;
ROM1[2670]<=26'd1953068; ROM2[2670]<=26'd11290068; ROM3[2670]<=26'd9753337; ROM4[2670]<=26'd23464568;
ROM1[2671]<=26'd1949658; ROM2[2671]<=26'd11289655; ROM3[2671]<=26'd9754623; ROM4[2671]<=26'd23463837;
ROM1[2672]<=26'd1950679; ROM2[2672]<=26'd11289416; ROM3[2672]<=26'd9752347; ROM4[2672]<=26'd23462424;
ROM1[2673]<=26'd1961028; ROM2[2673]<=26'd11291555; ROM3[2673]<=26'd9748380; ROM4[2673]<=26'd23463575;
ROM1[2674]<=26'd1971916; ROM2[2674]<=26'd11291055; ROM3[2674]<=26'd9740304; ROM4[2674]<=26'd23461523;
ROM1[2675]<=26'd1970991; ROM2[2675]<=26'd11289959; ROM3[2675]<=26'd9734273; ROM4[2675]<=26'd23459002;
ROM1[2676]<=26'd1966218; ROM2[2676]<=26'd11291839; ROM3[2676]<=26'd9736357; ROM4[2676]<=26'd23459253;
ROM1[2677]<=26'd1961615; ROM2[2677]<=26'd11294344; ROM3[2677]<=26'd9740950; ROM4[2677]<=26'd23460845;
ROM1[2678]<=26'd1956596; ROM2[2678]<=26'd11295527; ROM3[2678]<=26'd9742809; ROM4[2678]<=26'd23460330;
ROM1[2679]<=26'd1949340; ROM2[2679]<=26'd11292274; ROM3[2679]<=26'd9742474; ROM4[2679]<=26'd23456320;
ROM1[2680]<=26'd1946302; ROM2[2680]<=26'd11291016; ROM3[2680]<=26'd9738559; ROM4[2680]<=26'd23453990;
ROM1[2681]<=26'd1949999; ROM2[2681]<=26'd11291338; ROM3[2681]<=26'd9732835; ROM4[2681]<=26'd23451328;
ROM1[2682]<=26'd1959153; ROM2[2682]<=26'd11288522; ROM3[2682]<=26'd9721442; ROM4[2682]<=26'd23446501;
ROM1[2683]<=26'd1966072; ROM2[2683]<=26'd11290514; ROM3[2683]<=26'd9716220; ROM4[2683]<=26'd23446485;
ROM1[2684]<=26'd1962814; ROM2[2684]<=26'd11291598; ROM3[2684]<=26'd9717336; ROM4[2684]<=26'd23446563;
ROM1[2685]<=26'd1953425; ROM2[2685]<=26'd11287637; ROM3[2685]<=26'd9715810; ROM4[2685]<=26'd23443241;
ROM1[2686]<=26'd1950022; ROM2[2686]<=26'd11288861; ROM3[2686]<=26'd9722122; ROM4[2686]<=26'd23446072;
ROM1[2687]<=26'd1949822; ROM2[2687]<=26'd11293100; ROM3[2687]<=26'd9728674; ROM4[2687]<=26'd23451977;
ROM1[2688]<=26'd1946085; ROM2[2688]<=26'd11292249; ROM3[2688]<=26'd9728935; ROM4[2688]<=26'd23452719;
ROM1[2689]<=26'd1948568; ROM2[2689]<=26'd11292378; ROM3[2689]<=26'd9727739; ROM4[2689]<=26'd23452264;
ROM1[2690]<=26'd1958190; ROM2[2690]<=26'd11291116; ROM3[2690]<=26'd9722866; ROM4[2690]<=26'd23451309;
ROM1[2691]<=26'd1966415; ROM2[2691]<=26'd11288598; ROM3[2691]<=26'd9716778; ROM4[2691]<=26'd23448791;
ROM1[2692]<=26'd1961671; ROM2[2692]<=26'd11285625; ROM3[2692]<=26'd9715047; ROM4[2692]<=26'd23445405;
ROM1[2693]<=26'd1958703; ROM2[2693]<=26'd11289701; ROM3[2693]<=26'd9723722; ROM4[2693]<=26'd23450930;
ROM1[2694]<=26'd1955480; ROM2[2694]<=26'd11294821; ROM3[2694]<=26'd9732911; ROM4[2694]<=26'd23456353;
ROM1[2695]<=26'd1944661; ROM2[2695]<=26'd11288817; ROM3[2695]<=26'd9730906; ROM4[2695]<=26'd23451097;
ROM1[2696]<=26'd1940046; ROM2[2696]<=26'd11288010; ROM3[2696]<=26'd9733101; ROM4[2696]<=26'd23451675;
ROM1[2697]<=26'd1939789; ROM2[2697]<=26'd11287005; ROM3[2697]<=26'd9732427; ROM4[2697]<=26'd23451401;
ROM1[2698]<=26'd1943733; ROM2[2698]<=26'd11281841; ROM3[2698]<=26'd9724611; ROM4[2698]<=26'd23445843;
ROM1[2699]<=26'd1961193; ROM2[2699]<=26'd11289523; ROM3[2699]<=26'd9723096; ROM4[2699]<=26'd23450454;
ROM1[2700]<=26'd1975954; ROM2[2700]<=26'd11300461; ROM3[2700]<=26'd9730202; ROM4[2700]<=26'd23461433;
ROM1[2701]<=26'd1972698; ROM2[2701]<=26'd11300872; ROM3[2701]<=26'd9732495; ROM4[2701]<=26'd23462365;
ROM1[2702]<=26'd1956100; ROM2[2702]<=26'd11291955; ROM3[2702]<=26'd9727224; ROM4[2702]<=26'd23454396;
ROM1[2703]<=26'd1944873; ROM2[2703]<=26'd11286226; ROM3[2703]<=26'd9726683; ROM4[2703]<=26'd23450374;
ROM1[2704]<=26'd1933606; ROM2[2704]<=26'd11281565; ROM3[2704]<=26'd9727963; ROM4[2704]<=26'd23448235;
ROM1[2705]<=26'd1929519; ROM2[2705]<=26'd11280607; ROM3[2705]<=26'd9728017; ROM4[2705]<=26'd23447710;
ROM1[2706]<=26'd1941032; ROM2[2706]<=26'd11286408; ROM3[2706]<=26'd9730414; ROM4[2706]<=26'd23452982;
ROM1[2707]<=26'd1963410; ROM2[2707]<=26'd11296623; ROM3[2707]<=26'd9734155; ROM4[2707]<=26'd23462152;
ROM1[2708]<=26'd1968432; ROM2[2708]<=26'd11296134; ROM3[2708]<=26'd9728881; ROM4[2708]<=26'd23460263;
ROM1[2709]<=26'd1953773; ROM2[2709]<=26'd11284627; ROM3[2709]<=26'd9721780; ROM4[2709]<=26'd23449666;
ROM1[2710]<=26'd1946998; ROM2[2710]<=26'd11286255; ROM3[2710]<=26'd9727718; ROM4[2710]<=26'd23452167;
ROM1[2711]<=26'd1938851; ROM2[2711]<=26'd11285570; ROM3[2711]<=26'd9730014; ROM4[2711]<=26'd23450468;
ROM1[2712]<=26'd1928519; ROM2[2712]<=26'd11279933; ROM3[2712]<=26'd9728348; ROM4[2712]<=26'd23446219;
ROM1[2713]<=26'd1929543; ROM2[2713]<=26'd11283997; ROM3[2713]<=26'd9735429; ROM4[2713]<=26'd23451564;
ROM1[2714]<=26'd1941353; ROM2[2714]<=26'd11292876; ROM3[2714]<=26'd9742008; ROM4[2714]<=26'd23459128;
ROM1[2715]<=26'd1953384; ROM2[2715]<=26'd11294155; ROM3[2715]<=26'd9737345; ROM4[2715]<=26'd23460159;
ROM1[2716]<=26'd1960932; ROM2[2716]<=26'd11290778; ROM3[2716]<=26'd9728137; ROM4[2716]<=26'd23454656;
ROM1[2717]<=26'd1963828; ROM2[2717]<=26'd11295705; ROM3[2717]<=26'd9728406; ROM4[2717]<=26'd23458485;
ROM1[2718]<=26'd1957509; ROM2[2718]<=26'd11294575; ROM3[2718]<=26'd9729565; ROM4[2718]<=26'd23458279;
ROM1[2719]<=26'd1950791; ROM2[2719]<=26'd11291895; ROM3[2719]<=26'd9730778; ROM4[2719]<=26'd23456263;
ROM1[2720]<=26'd1945633; ROM2[2720]<=26'd11291782; ROM3[2720]<=26'd9734438; ROM4[2720]<=26'd23457336;
ROM1[2721]<=26'd1936605; ROM2[2721]<=26'd11288446; ROM3[2721]<=26'd9735777; ROM4[2721]<=26'd23456419;
ROM1[2722]<=26'd1935173; ROM2[2722]<=26'd11286783; ROM3[2722]<=26'd9732787; ROM4[2722]<=26'd23453523;
ROM1[2723]<=26'd1943190; ROM2[2723]<=26'd11287064; ROM3[2723]<=26'd9729008; ROM4[2723]<=26'd23452353;
ROM1[2724]<=26'd1959554; ROM2[2724]<=26'd11290789; ROM3[2724]<=26'd9726607; ROM4[2724]<=26'd23455467;
ROM1[2725]<=26'd1964205; ROM2[2725]<=26'd11290383; ROM3[2725]<=26'd9725750; ROM4[2725]<=26'd23456520;
ROM1[2726]<=26'd1958988; ROM2[2726]<=26'd11290557; ROM3[2726]<=26'd9731303; ROM4[2726]<=26'd23459512;
ROM1[2727]<=26'd1951547; ROM2[2727]<=26'd11292714; ROM3[2727]<=26'd9738876; ROM4[2727]<=26'd23461871;
ROM1[2728]<=26'd1948856; ROM2[2728]<=26'd11295010; ROM3[2728]<=26'd9744087; ROM4[2728]<=26'd23464560;
ROM1[2729]<=26'd1945474; ROM2[2729]<=26'd11296477; ROM3[2729]<=26'd9746609; ROM4[2729]<=26'd23463580;
ROM1[2730]<=26'd1938346; ROM2[2730]<=26'd11289985; ROM3[2730]<=26'd9740924; ROM4[2730]<=26'd23456426;
ROM1[2731]<=26'd1942136; ROM2[2731]<=26'd11287462; ROM3[2731]<=26'd9734627; ROM4[2731]<=26'd23454075;
ROM1[2732]<=26'd1959553; ROM2[2732]<=26'd11292904; ROM3[2732]<=26'd9731586; ROM4[2732]<=26'd23456035;
ROM1[2733]<=26'd1969808; ROM2[2733]<=26'd11295017; ROM3[2733]<=26'd9730024; ROM4[2733]<=26'd23458624;
ROM1[2734]<=26'd1966694; ROM2[2734]<=26'd11296754; ROM3[2734]<=26'd9731749; ROM4[2734]<=26'd23460671;
ROM1[2735]<=26'd1963366; ROM2[2735]<=26'd11297703; ROM3[2735]<=26'd9737511; ROM4[2735]<=26'd23463005;
ROM1[2736]<=26'd1956152; ROM2[2736]<=26'd11294145; ROM3[2736]<=26'd9741471; ROM4[2736]<=26'd23462184;
ROM1[2737]<=26'd1949066; ROM2[2737]<=26'd11293558; ROM3[2737]<=26'd9742748; ROM4[2737]<=26'd23460624;
ROM1[2738]<=26'd1946041; ROM2[2738]<=26'd11295116; ROM3[2738]<=26'd9744317; ROM4[2738]<=26'd23461598;
ROM1[2739]<=26'd1946549; ROM2[2739]<=26'd11293873; ROM3[2739]<=26'd9742590; ROM4[2739]<=26'd23460680;
ROM1[2740]<=26'd1956208; ROM2[2740]<=26'd11295988; ROM3[2740]<=26'd9738892; ROM4[2740]<=26'd23461205;
ROM1[2741]<=26'd1970364; ROM2[2741]<=26'd11298919; ROM3[2741]<=26'd9736791; ROM4[2741]<=26'd23463781;
ROM1[2742]<=26'd1970833; ROM2[2742]<=26'd11298859; ROM3[2742]<=26'd9736495; ROM4[2742]<=26'd23464022;
ROM1[2743]<=26'd1962341; ROM2[2743]<=26'd11297283; ROM3[2743]<=26'd9736598; ROM4[2743]<=26'd23463624;
ROM1[2744]<=26'd1957621; ROM2[2744]<=26'd11297925; ROM3[2744]<=26'd9740725; ROM4[2744]<=26'd23466154;
ROM1[2745]<=26'd1953362; ROM2[2745]<=26'd11299996; ROM3[2745]<=26'd9745827; ROM4[2745]<=26'd23469240;
ROM1[2746]<=26'd1951278; ROM2[2746]<=26'd11303393; ROM3[2746]<=26'd9752229; ROM4[2746]<=26'd23474640;
ROM1[2747]<=26'd1957049; ROM2[2747]<=26'd11307162; ROM3[2747]<=26'd9757250; ROM4[2747]<=26'd23477916;
ROM1[2748]<=26'd1961704; ROM2[2748]<=26'd11303866; ROM3[2748]<=26'd9752483; ROM4[2748]<=26'd23474858;
ROM1[2749]<=26'd1971684; ROM2[2749]<=26'd11301336; ROM3[2749]<=26'd9746040; ROM4[2749]<=26'd23474346;
ROM1[2750]<=26'd1976394; ROM2[2750]<=26'd11302692; ROM3[2750]<=26'd9748478; ROM4[2750]<=26'd23478517;
ROM1[2751]<=26'd1973038; ROM2[2751]<=26'd11309017; ROM3[2751]<=26'd9754855; ROM4[2751]<=26'd23485184;
ROM1[2752]<=26'd1968006; ROM2[2752]<=26'd11311976; ROM3[2752]<=26'd9756455; ROM4[2752]<=26'd23486448;
ROM1[2753]<=26'd1961656; ROM2[2753]<=26'd11308303; ROM3[2753]<=26'd9752664; ROM4[2753]<=26'd23481483;
ROM1[2754]<=26'd1957560; ROM2[2754]<=26'd11308878; ROM3[2754]<=26'd9754682; ROM4[2754]<=26'd23480778;
ROM1[2755]<=26'd1951081; ROM2[2755]<=26'd11301894; ROM3[2755]<=26'd9750584; ROM4[2755]<=26'd23476176;
ROM1[2756]<=26'd1949878; ROM2[2756]<=26'd11296157; ROM3[2756]<=26'd9741712; ROM4[2756]<=26'd23470006;
ROM1[2757]<=26'd1961725; ROM2[2757]<=26'd11300263; ROM3[2757]<=26'd9736661; ROM4[2757]<=26'd23470585;
ROM1[2758]<=26'd1971904; ROM2[2758]<=26'd11302092; ROM3[2758]<=26'd9733457; ROM4[2758]<=26'd23470735;
ROM1[2759]<=26'd1977045; ROM2[2759]<=26'd11309826; ROM3[2759]<=26'd9740870; ROM4[2759]<=26'd23476371;
ROM1[2760]<=26'd1968943; ROM2[2760]<=26'd11309707; ROM3[2760]<=26'd9744328; ROM4[2760]<=26'd23476627;
ROM1[2761]<=26'd1953534; ROM2[2761]<=26'd11300497; ROM3[2761]<=26'd9740180; ROM4[2761]<=26'd23469365;
ROM1[2762]<=26'd1941943; ROM2[2762]<=26'd11293562; ROM3[2762]<=26'd9736249; ROM4[2762]<=26'd23464536;
ROM1[2763]<=26'd1934311; ROM2[2763]<=26'd11289168; ROM3[2763]<=26'd9732976; ROM4[2763]<=26'd23459570;
ROM1[2764]<=26'd1937981; ROM2[2764]<=26'd11290787; ROM3[2764]<=26'd9731464; ROM4[2764]<=26'd23458799;
ROM1[2765]<=26'd1952630; ROM2[2765]<=26'd11294919; ROM3[2765]<=26'd9730558; ROM4[2765]<=26'd23461667;
ROM1[2766]<=26'd1962185; ROM2[2766]<=26'd11294037; ROM3[2766]<=26'd9723795; ROM4[2766]<=26'd23458587;
ROM1[2767]<=26'd1954838; ROM2[2767]<=26'd11288338; ROM3[2767]<=26'd9717169; ROM4[2767]<=26'd23451667;
ROM1[2768]<=26'd1951275; ROM2[2768]<=26'd11290196; ROM3[2768]<=26'd9721832; ROM4[2768]<=26'd23455443;
ROM1[2769]<=26'd1948345; ROM2[2769]<=26'd11292998; ROM3[2769]<=26'd9729612; ROM4[2769]<=26'd23459756;
ROM1[2770]<=26'd1938860; ROM2[2770]<=26'd11291082; ROM3[2770]<=26'd9731990; ROM4[2770]<=26'd23457432;
ROM1[2771]<=26'd1930390; ROM2[2771]<=26'd11286390; ROM3[2771]<=26'd9732455; ROM4[2771]<=26'd23454664;
ROM1[2772]<=26'd1930504; ROM2[2772]<=26'd11285385; ROM3[2772]<=26'd9733000; ROM4[2772]<=26'd23453483;
ROM1[2773]<=26'd1939905; ROM2[2773]<=26'd11287864; ROM3[2773]<=26'd9728692; ROM4[2773]<=26'd23453122;
ROM1[2774]<=26'd1951466; ROM2[2774]<=26'd11286837; ROM3[2774]<=26'd9723173; ROM4[2774]<=26'd23451787;
ROM1[2775]<=26'd1954724; ROM2[2775]<=26'd11287468; ROM3[2775]<=26'd9722188; ROM4[2775]<=26'd23451564;
ROM1[2776]<=26'd1954452; ROM2[2776]<=26'd11291195; ROM3[2776]<=26'd9728009; ROM4[2776]<=26'd23455442;
ROM1[2777]<=26'd1949693; ROM2[2777]<=26'd11292489; ROM3[2777]<=26'd9734164; ROM4[2777]<=26'd23456488;
ROM1[2778]<=26'd1944730; ROM2[2778]<=26'd11291938; ROM3[2778]<=26'd9735664; ROM4[2778]<=26'd23456340;
ROM1[2779]<=26'd1940086; ROM2[2779]<=26'd11290241; ROM3[2779]<=26'd9739078; ROM4[2779]<=26'd23457166;
ROM1[2780]<=26'd1936392; ROM2[2780]<=26'd11287559; ROM3[2780]<=26'd9739150; ROM4[2780]<=26'd23455891;
ROM1[2781]<=26'd1940402; ROM2[2781]<=26'd11287932; ROM3[2781]<=26'd9737415; ROM4[2781]<=26'd23455697;
ROM1[2782]<=26'd1955371; ROM2[2782]<=26'd11292070; ROM3[2782]<=26'd9734758; ROM4[2782]<=26'd23458130;
ROM1[2783]<=26'd1969483; ROM2[2783]<=26'd11299307; ROM3[2783]<=26'd9735323; ROM4[2783]<=26'd23463541;
ROM1[2784]<=26'd1974088; ROM2[2784]<=26'd11306078; ROM3[2784]<=26'd9742886; ROM4[2784]<=26'd23468856;
ROM1[2785]<=26'd1964013; ROM2[2785]<=26'd11300081; ROM3[2785]<=26'd9741283; ROM4[2785]<=26'd23463955;
ROM1[2786]<=26'd1955152; ROM2[2786]<=26'd11293685; ROM3[2786]<=26'd9740255; ROM4[2786]<=26'd23459575;
ROM1[2787]<=26'd1953191; ROM2[2787]<=26'd11295778; ROM3[2787]<=26'd9745901; ROM4[2787]<=26'd23463400;
ROM1[2788]<=26'd1947536; ROM2[2788]<=26'd11293992; ROM3[2788]<=26'd9745234; ROM4[2788]<=26'd23462245;
ROM1[2789]<=26'd1955138; ROM2[2789]<=26'd11297613; ROM3[2789]<=26'd9748312; ROM4[2789]<=26'd23467413;
ROM1[2790]<=26'd1978823; ROM2[2790]<=26'd11311306; ROM3[2790]<=26'd9758285; ROM4[2790]<=26'd23480781;
ROM1[2791]<=26'd1989113; ROM2[2791]<=26'd11312816; ROM3[2791]<=26'd9752198; ROM4[2791]<=26'd23479810;
ROM1[2792]<=26'd1979547; ROM2[2792]<=26'd11302575; ROM3[2792]<=26'd9740492; ROM4[2792]<=26'd23470192;
ROM1[2793]<=26'd1969464; ROM2[2793]<=26'd11299255; ROM3[2793]<=26'd9740505; ROM4[2793]<=26'd23467486;
ROM1[2794]<=26'd1959294; ROM2[2794]<=26'd11296715; ROM3[2794]<=26'd9740179; ROM4[2794]<=26'd23464739;
ROM1[2795]<=26'd1953894; ROM2[2795]<=26'd11294681; ROM3[2795]<=26'd9742183; ROM4[2795]<=26'd23465680;
ROM1[2796]<=26'd1952108; ROM2[2796]<=26'd11299074; ROM3[2796]<=26'd9749172; ROM4[2796]<=26'd23469946;
ROM1[2797]<=26'd1955476; ROM2[2797]<=26'd11302470; ROM3[2797]<=26'd9749910; ROM4[2797]<=26'd23470538;
ROM1[2798]<=26'd1962729; ROM2[2798]<=26'd11303082; ROM3[2798]<=26'd9742406; ROM4[2798]<=26'd23466802;
ROM1[2799]<=26'd1972264; ROM2[2799]<=26'd11301149; ROM3[2799]<=26'd9735045; ROM4[2799]<=26'd23463295;
ROM1[2800]<=26'd1974661; ROM2[2800]<=26'd11300454; ROM3[2800]<=26'd9736436; ROM4[2800]<=26'd23466439;
ROM1[2801]<=26'd1972356; ROM2[2801]<=26'd11303739; ROM3[2801]<=26'd9745234; ROM4[2801]<=26'd23472118;
ROM1[2802]<=26'd1967171; ROM2[2802]<=26'd11303952; ROM3[2802]<=26'd9750927; ROM4[2802]<=26'd23473296;
ROM1[2803]<=26'd1965576; ROM2[2803]<=26'd11306686; ROM3[2803]<=26'd9758477; ROM4[2803]<=26'd23477475;
ROM1[2804]<=26'd1963605; ROM2[2804]<=26'd11308388; ROM3[2804]<=26'd9765303; ROM4[2804]<=26'd23481054;
ROM1[2805]<=26'd1956571; ROM2[2805]<=26'd11303149; ROM3[2805]<=26'd9761501; ROM4[2805]<=26'd23476371;
ROM1[2806]<=26'd1958414; ROM2[2806]<=26'd11301296; ROM3[2806]<=26'd9756719; ROM4[2806]<=26'd23473149;
ROM1[2807]<=26'd1968372; ROM2[2807]<=26'd11300933; ROM3[2807]<=26'd9746987; ROM4[2807]<=26'd23469774;
ROM1[2808]<=26'd1974244; ROM2[2808]<=26'd11299778; ROM3[2808]<=26'd9741391; ROM4[2808]<=26'd23467609;
ROM1[2809]<=26'd1975372; ROM2[2809]<=26'd11303274; ROM3[2809]<=26'd9746484; ROM4[2809]<=26'd23471739;
ROM1[2810]<=26'd1965517; ROM2[2810]<=26'd11300810; ROM3[2810]<=26'd9748333; ROM4[2810]<=26'd23472637;
ROM1[2811]<=26'd1956221; ROM2[2811]<=26'd11299441; ROM3[2811]<=26'd9750436; ROM4[2811]<=26'd23471445;
ROM1[2812]<=26'd1952728; ROM2[2812]<=26'd11300961; ROM3[2812]<=26'd9754152; ROM4[2812]<=26'd23473783;
ROM1[2813]<=26'd1949533; ROM2[2813]<=26'd11300714; ROM3[2813]<=26'd9756315; ROM4[2813]<=26'd23474165;
ROM1[2814]<=26'd1955586; ROM2[2814]<=26'd11303915; ROM3[2814]<=26'd9758174; ROM4[2814]<=26'd23475900;
ROM1[2815]<=26'd1965840; ROM2[2815]<=26'd11303743; ROM3[2815]<=26'd9753541; ROM4[2815]<=26'd23475823;
ROM1[2816]<=26'd1974944; ROM2[2816]<=26'd11302594; ROM3[2816]<=26'd9745699; ROM4[2816]<=26'd23473167;
ROM1[2817]<=26'd1974371; ROM2[2817]<=26'd11303830; ROM3[2817]<=26'd9744455; ROM4[2817]<=26'd23473200;
ROM1[2818]<=26'd1967577; ROM2[2818]<=26'd11302637; ROM3[2818]<=26'd9748652; ROM4[2818]<=26'd23472858;
ROM1[2819]<=26'd1962918; ROM2[2819]<=26'd11304297; ROM3[2819]<=26'd9754282; ROM4[2819]<=26'd23476811;
ROM1[2820]<=26'd1961413; ROM2[2820]<=26'd11310259; ROM3[2820]<=26'd9759556; ROM4[2820]<=26'd23480862;
ROM1[2821]<=26'd1952493; ROM2[2821]<=26'd11306020; ROM3[2821]<=26'd9756444; ROM4[2821]<=26'd23475806;
ROM1[2822]<=26'd1952001; ROM2[2822]<=26'd11302365; ROM3[2822]<=26'd9752697; ROM4[2822]<=26'd23473016;
ROM1[2823]<=26'd1962271; ROM2[2823]<=26'd11303251; ROM3[2823]<=26'd9750924; ROM4[2823]<=26'd23472986;
ROM1[2824]<=26'd1971710; ROM2[2824]<=26'd11301745; ROM3[2824]<=26'd9745293; ROM4[2824]<=26'd23471326;
ROM1[2825]<=26'd1975887; ROM2[2825]<=26'd11301351; ROM3[2825]<=26'd9745288; ROM4[2825]<=26'd23473073;
ROM1[2826]<=26'd1972200; ROM2[2826]<=26'd11303154; ROM3[2826]<=26'd9748207; ROM4[2826]<=26'd23474970;
ROM1[2827]<=26'd1967081; ROM2[2827]<=26'd11303866; ROM3[2827]<=26'd9751481; ROM4[2827]<=26'd23474192;
ROM1[2828]<=26'd1963896; ROM2[2828]<=26'd11302343; ROM3[2828]<=26'd9755002; ROM4[2828]<=26'd23473481;
ROM1[2829]<=26'd1958100; ROM2[2829]<=26'd11302887; ROM3[2829]<=26'd9757783; ROM4[2829]<=26'd23474097;
ROM1[2830]<=26'd1954004; ROM2[2830]<=26'd11302000; ROM3[2830]<=26'd9754931; ROM4[2830]<=26'd23473666;
ROM1[2831]<=26'd1957430; ROM2[2831]<=26'd11298806; ROM3[2831]<=26'd9748790; ROM4[2831]<=26'd23469365;
ROM1[2832]<=26'd1968202; ROM2[2832]<=26'd11296687; ROM3[2832]<=26'd9740022; ROM4[2832]<=26'd23465349;
ROM1[2833]<=26'd1976113; ROM2[2833]<=26'd11298353; ROM3[2833]<=26'd9736613; ROM4[2833]<=26'd23466966;
ROM1[2834]<=26'd1973012; ROM2[2834]<=26'd11300621; ROM3[2834]<=26'd9741620; ROM4[2834]<=26'd23467958;
ROM1[2835]<=26'd1963482; ROM2[2835]<=26'd11300755; ROM3[2835]<=26'd9743356; ROM4[2835]<=26'd23467473;
ROM1[2836]<=26'd1955652; ROM2[2836]<=26'd11299273; ROM3[2836]<=26'd9745111; ROM4[2836]<=26'd23466834;
ROM1[2837]<=26'd1945303; ROM2[2837]<=26'd11291590; ROM3[2837]<=26'd9742953; ROM4[2837]<=26'd23459615;
ROM1[2838]<=26'd1937532; ROM2[2838]<=26'd11287884; ROM3[2838]<=26'd9739633; ROM4[2838]<=26'd23454858;
ROM1[2839]<=26'd1937233; ROM2[2839]<=26'd11285483; ROM3[2839]<=26'd9736201; ROM4[2839]<=26'd23451525;
ROM1[2840]<=26'd1948084; ROM2[2840]<=26'd11287432; ROM3[2840]<=26'd9730866; ROM4[2840]<=26'd23449261;
ROM1[2841]<=26'd1964083; ROM2[2841]<=26'd11296140; ROM3[2841]<=26'd9730781; ROM4[2841]<=26'd23454065;
ROM1[2842]<=26'd1971805; ROM2[2842]<=26'd11302512; ROM3[2842]<=26'd9736451; ROM4[2842]<=26'd23459480;
ROM1[2843]<=26'd1966025; ROM2[2843]<=26'd11304613; ROM3[2843]<=26'd9740662; ROM4[2843]<=26'd23460903;
ROM1[2844]<=26'd1948071; ROM2[2844]<=26'd11296121; ROM3[2844]<=26'd9736858; ROM4[2844]<=26'd23454240;
ROM1[2845]<=26'd1937954; ROM2[2845]<=26'd11289986; ROM3[2845]<=26'd9736025; ROM4[2845]<=26'd23450097;
ROM1[2846]<=26'd1929801; ROM2[2846]<=26'd11287219; ROM3[2846]<=26'd9735647; ROM4[2846]<=26'd23447352;
ROM1[2847]<=26'd1931164; ROM2[2847]<=26'd11286115; ROM3[2847]<=26'd9734070; ROM4[2847]<=26'd23445843;
ROM1[2848]<=26'd1948271; ROM2[2848]<=26'd11294391; ROM3[2848]<=26'd9738287; ROM4[2848]<=26'd23452182;
ROM1[2849]<=26'd1963940; ROM2[2849]<=26'd11299329; ROM3[2849]<=26'd9737019; ROM4[2849]<=26'd23455457;
ROM1[2850]<=26'd1961913; ROM2[2850]<=26'd11293250; ROM3[2850]<=26'd9727965; ROM4[2850]<=26'd23451017;
ROM1[2851]<=26'd1953388; ROM2[2851]<=26'd11289079; ROM3[2851]<=26'd9726758; ROM4[2851]<=26'd23449168;
ROM1[2852]<=26'd1946258; ROM2[2852]<=26'd11287565; ROM3[2852]<=26'd9730368; ROM4[2852]<=26'd23450240;
ROM1[2853]<=26'd1940975; ROM2[2853]<=26'd11287305; ROM3[2853]<=26'd9731964; ROM4[2853]<=26'd23448771;
ROM1[2854]<=26'd1937221; ROM2[2854]<=26'd11289387; ROM3[2854]<=26'd9738727; ROM4[2854]<=26'd23453221;
ROM1[2855]<=26'd1935541; ROM2[2855]<=26'd11289399; ROM3[2855]<=26'd9742660; ROM4[2855]<=26'd23455999;
ROM1[2856]<=26'd1947151; ROM2[2856]<=26'd11295126; ROM3[2856]<=26'd9745522; ROM4[2856]<=26'd23460688;
ROM1[2857]<=26'd1969500; ROM2[2857]<=26'd11305859; ROM3[2857]<=26'd9748394; ROM4[2857]<=26'd23470441;
ROM1[2858]<=26'd1976560; ROM2[2858]<=26'd11306474; ROM3[2858]<=26'd9744343; ROM4[2858]<=26'd23468994;
ROM1[2859]<=26'd1969069; ROM2[2859]<=26'd11301941; ROM3[2859]<=26'd9741790; ROM4[2859]<=26'd23465492;
ROM1[2860]<=26'd1960563; ROM2[2860]<=26'd11299723; ROM3[2860]<=26'd9743180; ROM4[2860]<=26'd23464067;
ROM1[2861]<=26'd1953778; ROM2[2861]<=26'd11297328; ROM3[2861]<=26'd9744948; ROM4[2861]<=26'd23462669;
ROM1[2862]<=26'd1950127; ROM2[2862]<=26'd11298237; ROM3[2862]<=26'd9749742; ROM4[2862]<=26'd23464648;
ROM1[2863]<=26'd1949572; ROM2[2863]<=26'd11301628; ROM3[2863]<=26'd9753456; ROM4[2863]<=26'd23465925;
ROM1[2864]<=26'd1953540; ROM2[2864]<=26'd11303505; ROM3[2864]<=26'd9752442; ROM4[2864]<=26'd23466575;
ROM1[2865]<=26'd1960607; ROM2[2865]<=26'd11301836; ROM3[2865]<=26'd9745338; ROM4[2865]<=26'd23463132;
ROM1[2866]<=26'd1972416; ROM2[2866]<=26'd11304084; ROM3[2866]<=26'd9742995; ROM4[2866]<=26'd23464648;
ROM1[2867]<=26'd1980852; ROM2[2867]<=26'd11312411; ROM3[2867]<=26'd9752013; ROM4[2867]<=26'd23473843;
ROM1[2868]<=26'd1970754; ROM2[2868]<=26'd11309642; ROM3[2868]<=26'd9752997; ROM4[2868]<=26'd23471366;
ROM1[2869]<=26'd1958422; ROM2[2869]<=26'd11302316; ROM3[2869]<=26'd9750177; ROM4[2869]<=26'd23466222;
ROM1[2870]<=26'd1956951; ROM2[2870]<=26'd11302940; ROM3[2870]<=26'd9755361; ROM4[2870]<=26'd23468952;
ROM1[2871]<=26'd1962296; ROM2[2871]<=26'd11311956; ROM3[2871]<=26'd9767978; ROM4[2871]<=26'd23478153;
ROM1[2872]<=26'd1967069; ROM2[2872]<=26'd11313613; ROM3[2872]<=26'd9770802; ROM4[2872]<=26'd23482180;
ROM1[2873]<=26'd1972592; ROM2[2873]<=26'd11310030; ROM3[2873]<=26'd9764297; ROM4[2873]<=26'd23479702;
ROM1[2874]<=26'd1985827; ROM2[2874]<=26'd11312103; ROM3[2874]<=26'd9759153; ROM4[2874]<=26'd23479819;
ROM1[2875]<=26'd1983968; ROM2[2875]<=26'd11308687; ROM3[2875]<=26'd9752769; ROM4[2875]<=26'd23476249;
ROM1[2876]<=26'd1973056; ROM2[2876]<=26'd11302380; ROM3[2876]<=26'd9748766; ROM4[2876]<=26'd23470496;
ROM1[2877]<=26'd1967820; ROM2[2877]<=26'd11300601; ROM3[2877]<=26'd9751600; ROM4[2877]<=26'd23469756;
ROM1[2878]<=26'd1962115; ROM2[2878]<=26'd11301320; ROM3[2878]<=26'd9754940; ROM4[2878]<=26'd23471299;
ROM1[2879]<=26'd1950323; ROM2[2879]<=26'd11297257; ROM3[2879]<=26'd9753076; ROM4[2879]<=26'd23466667;
ROM1[2880]<=26'd1949867; ROM2[2880]<=26'd11296839; ROM3[2880]<=26'd9753321; ROM4[2880]<=26'd23466907;
ROM1[2881]<=26'd1962562; ROM2[2881]<=26'd11302288; ROM3[2881]<=26'd9755732; ROM4[2881]<=26'd23473340;
ROM1[2882]<=26'd1981024; ROM2[2882]<=26'd11305445; ROM3[2882]<=26'd9752683; ROM4[2882]<=26'd23474800;
ROM1[2883]<=26'd1984716; ROM2[2883]<=26'd11300798; ROM3[2883]<=26'd9742540; ROM4[2883]<=26'd23468878;
ROM1[2884]<=26'd1979740; ROM2[2884]<=26'd11302629; ROM3[2884]<=26'd9743107; ROM4[2884]<=26'd23470478;
ROM1[2885]<=26'd1975929; ROM2[2885]<=26'd11307441; ROM3[2885]<=26'd9749819; ROM4[2885]<=26'd23474379;
ROM1[2886]<=26'd1973065; ROM2[2886]<=26'd11308323; ROM3[2886]<=26'd9753639; ROM4[2886]<=26'd23475619;
ROM1[2887]<=26'd1976884; ROM2[2887]<=26'd11314281; ROM3[2887]<=26'd9764562; ROM4[2887]<=26'd23482539;
ROM1[2888]<=26'd1977756; ROM2[2888]<=26'd11318694; ROM3[2888]<=26'd9771994; ROM4[2888]<=26'd23486949;
ROM1[2889]<=26'd1977090; ROM2[2889]<=26'd11316376; ROM3[2889]<=26'd9767581; ROM4[2889]<=26'd23483365;
ROM1[2890]<=26'd1992984; ROM2[2890]<=26'd11315275; ROM3[2890]<=26'd9759112; ROM4[2890]<=26'd23479523;
ROM1[2891]<=26'd2009667; ROM2[2891]<=26'd11317475; ROM3[2891]<=26'd9751323; ROM4[2891]<=26'd23478942;
ROM1[2892]<=26'd2011389; ROM2[2892]<=26'd11317014; ROM3[2892]<=26'd9749169; ROM4[2892]<=26'd23477288;
ROM1[2893]<=26'd2011481; ROM2[2893]<=26'd11318426; ROM3[2893]<=26'd9756372; ROM4[2893]<=26'd23480744;
ROM1[2894]<=26'd2008526; ROM2[2894]<=26'd11318748; ROM3[2894]<=26'd9763469; ROM4[2894]<=26'd23483171;
ROM1[2895]<=26'd2007298; ROM2[2895]<=26'd11319088; ROM3[2895]<=26'd9767911; ROM4[2895]<=26'd23485302;
ROM1[2896]<=26'd2011836; ROM2[2896]<=26'd11322934; ROM3[2896]<=26'd9774961; ROM4[2896]<=26'd23491056;
ROM1[2897]<=26'd2023610; ROM2[2897]<=26'd11328665; ROM3[2897]<=26'd9776593; ROM4[2897]<=26'd23495717;
ROM1[2898]<=26'd2038234; ROM2[2898]<=26'd11332574; ROM3[2898]<=26'd9772799; ROM4[2898]<=26'd23497738;
ROM1[2899]<=26'd2058713; ROM2[2899]<=26'd11336112; ROM3[2899]<=26'd9766988; ROM4[2899]<=26'd23498371;
ROM1[2900]<=26'd2074186; ROM2[2900]<=26'd11342570; ROM3[2900]<=26'd9766690; ROM4[2900]<=26'd23501261;
ROM1[2901]<=26'd2085154; ROM2[2901]<=26'd11354499; ROM3[2901]<=26'd9776957; ROM4[2901]<=26'd23511074;
ROM1[2902]<=26'd2086589; ROM2[2902]<=26'd11358600; ROM3[2902]<=26'd9784513; ROM4[2902]<=26'd23517064;
ROM1[2903]<=26'd2085718; ROM2[2903]<=26'd11357030; ROM3[2903]<=26'd9786198; ROM4[2903]<=26'd23516897;
ROM1[2904]<=26'd2081072; ROM2[2904]<=26'd11355404; ROM3[2904]<=26'd9783111; ROM4[2904]<=26'd23513108;
ROM1[2905]<=26'd2077669; ROM2[2905]<=26'd11351329; ROM3[2905]<=26'd9774856; ROM4[2905]<=26'd23506341;
ROM1[2906]<=26'd2082886; ROM2[2906]<=26'd11349374; ROM3[2906]<=26'd9766653; ROM4[2906]<=26'd23501169;
ROM1[2907]<=26'd2099584; ROM2[2907]<=26'd11351426; ROM3[2907]<=26'd9760056; ROM4[2907]<=26'd23500862;
ROM1[2908]<=26'd2112135; ROM2[2908]<=26'd11351504; ROM3[2908]<=26'd9758614; ROM4[2908]<=26'd23501312;
ROM1[2909]<=26'd2109761; ROM2[2909]<=26'd11348186; ROM3[2909]<=26'd9759131; ROM4[2909]<=26'd23499003;
ROM1[2910]<=26'd2104241; ROM2[2910]<=26'd11348375; ROM3[2910]<=26'd9761273; ROM4[2910]<=26'd23500203;
ROM1[2911]<=26'd2102172; ROM2[2911]<=26'd11350108; ROM3[2911]<=26'd9763774; ROM4[2911]<=26'd23500911;
ROM1[2912]<=26'd2102519; ROM2[2912]<=26'd11351658; ROM3[2912]<=26'd9764098; ROM4[2912]<=26'd23501500;
ROM1[2913]<=26'd2107405; ROM2[2913]<=26'd11358290; ROM3[2913]<=26'd9767893; ROM4[2913]<=26'd23505903;
ROM1[2914]<=26'd2120152; ROM2[2914]<=26'd11366221; ROM3[2914]<=26'd9770979; ROM4[2914]<=26'd23510077;
ROM1[2915]<=26'd2139485; ROM2[2915]<=26'd11373878; ROM3[2915]<=26'd9770761; ROM4[2915]<=26'd23515310;
ROM1[2916]<=26'd2155426; ROM2[2916]<=26'd11376884; ROM3[2916]<=26'd9768909; ROM4[2916]<=26'd23517141;
ROM1[2917]<=26'd2153537; ROM2[2917]<=26'd11371702; ROM3[2917]<=26'd9765336; ROM4[2917]<=26'd23513723;
ROM1[2918]<=26'd2147788; ROM2[2918]<=26'd11373033; ROM3[2918]<=26'd9767540; ROM4[2918]<=26'd23513181;
ROM1[2919]<=26'd2148520; ROM2[2919]<=26'd11377698; ROM3[2919]<=26'd9774810; ROM4[2919]<=26'd23516457;
ROM1[2920]<=26'd2146258; ROM2[2920]<=26'd11373487; ROM3[2920]<=26'd9773505; ROM4[2920]<=26'd23514093;
ROM1[2921]<=26'd2140220; ROM2[2921]<=26'd11365991; ROM3[2921]<=26'd9770044; ROM4[2921]<=26'd23508134;
ROM1[2922]<=26'd2148660; ROM2[2922]<=26'd11367935; ROM3[2922]<=26'd9771309; ROM4[2922]<=26'd23510218;
ROM1[2923]<=26'd2161612; ROM2[2923]<=26'd11370685; ROM3[2923]<=26'd9768207; ROM4[2923]<=26'd23513246;
ROM1[2924]<=26'd2176588; ROM2[2924]<=26'd11374365; ROM3[2924]<=26'd9763552; ROM4[2924]<=26'd23515571;
ROM1[2925]<=26'd2182882; ROM2[2925]<=26'd11378269; ROM3[2925]<=26'd9763558; ROM4[2925]<=26'd23518264;
ROM1[2926]<=26'd2181334; ROM2[2926]<=26'd11377067; ROM3[2926]<=26'd9764131; ROM4[2926]<=26'd23519504;
ROM1[2927]<=26'd2178208; ROM2[2927]<=26'd11374838; ROM3[2927]<=26'd9767509; ROM4[2927]<=26'd23520326;
ROM1[2928]<=26'd2177196; ROM2[2928]<=26'd11378918; ROM3[2928]<=26'd9773933; ROM4[2928]<=26'd23525360;
ROM1[2929]<=26'd2183298; ROM2[2929]<=26'd11391816; ROM3[2929]<=26'd9785625; ROM4[2929]<=26'd23535411;
ROM1[2930]<=26'd2190512; ROM2[2930]<=26'd11397208; ROM3[2930]<=26'd9791731; ROM4[2930]<=26'd23540563;
ROM1[2931]<=26'd2188535; ROM2[2931]<=26'd11389872; ROM3[2931]<=26'd9781169; ROM4[2931]<=26'd23534077;
ROM1[2932]<=26'd2197161; ROM2[2932]<=26'd11385968; ROM3[2932]<=26'd9772124; ROM4[2932]<=26'd23527928;
ROM1[2933]<=26'd2209818; ROM2[2933]<=26'd11388968; ROM3[2933]<=26'd9773082; ROM4[2933]<=26'd23531337;
ROM1[2934]<=26'd2204542; ROM2[2934]<=26'd11388998; ROM3[2934]<=26'd9773978; ROM4[2934]<=26'd23531450;
ROM1[2935]<=26'd2198324; ROM2[2935]<=26'd11389405; ROM3[2935]<=26'd9778782; ROM4[2935]<=26'd23532022;
ROM1[2936]<=26'd2200875; ROM2[2936]<=26'd11395405; ROM3[2936]<=26'd9790366; ROM4[2936]<=26'd23540350;
ROM1[2937]<=26'd2193517; ROM2[2937]<=26'd11392836; ROM3[2937]<=26'd9792515; ROM4[2937]<=26'd23539774;
ROM1[2938]<=26'd2185034; ROM2[2938]<=26'd11387349; ROM3[2938]<=26'd9789511; ROM4[2938]<=26'd23534936;
ROM1[2939]<=26'd2190218; ROM2[2939]<=26'd11387707; ROM3[2939]<=26'd9790699; ROM4[2939]<=26'd23536514;
ROM1[2940]<=26'd2202777; ROM2[2940]<=26'd11388871; ROM3[2940]<=26'd9787644; ROM4[2940]<=26'd23537867;
ROM1[2941]<=26'd2215983; ROM2[2941]<=26'd11391554; ROM3[2941]<=26'd9784152; ROM4[2941]<=26'd23538426;
ROM1[2942]<=26'd2216570; ROM2[2942]<=26'd11395178; ROM3[2942]<=26'd9787000; ROM4[2942]<=26'd23540464;
ROM1[2943]<=26'd2213209; ROM2[2943]<=26'd11399491; ROM3[2943]<=26'd9794332; ROM4[2943]<=26'd23544923;
ROM1[2944]<=26'd2205284; ROM2[2944]<=26'd11398994; ROM3[2944]<=26'd9797375; ROM4[2944]<=26'd23545013;
ROM1[2945]<=26'd2191338; ROM2[2945]<=26'd11390325; ROM3[2945]<=26'd9793648; ROM4[2945]<=26'd23538770;
ROM1[2946]<=26'd2180545; ROM2[2946]<=26'd11383438; ROM3[2946]<=26'd9790675; ROM4[2946]<=26'd23535267;
ROM1[2947]<=26'd2177976; ROM2[2947]<=26'd11381894; ROM3[2947]<=26'd9787591; ROM4[2947]<=26'd23533289;
ROM1[2948]<=26'd2182747; ROM2[2948]<=26'd11381542; ROM3[2948]<=26'd9783791; ROM4[2948]<=26'd23531581;
ROM1[2949]<=26'd2195955; ROM2[2949]<=26'd11383071; ROM3[2949]<=26'd9779296; ROM4[2949]<=26'd23532805;
ROM1[2950]<=26'd2197723; ROM2[2950]<=26'd11382162; ROM3[2950]<=26'd9777538; ROM4[2950]<=26'd23531440;
ROM1[2951]<=26'd2188512; ROM2[2951]<=26'd11378243; ROM3[2951]<=26'd9778466; ROM4[2951]<=26'd23527693;
ROM1[2952]<=26'd2182384; ROM2[2952]<=26'd11378375; ROM3[2952]<=26'd9783684; ROM4[2952]<=26'd23529497;
ROM1[2953]<=26'd2179370; ROM2[2953]<=26'd11381420; ROM3[2953]<=26'd9789939; ROM4[2953]<=26'd23535154;
ROM1[2954]<=26'd2169857; ROM2[2954]<=26'd11379376; ROM3[2954]<=26'd9792768; ROM4[2954]<=26'd23536941;
ROM1[2955]<=26'd2161654; ROM2[2955]<=26'd11376645; ROM3[2955]<=26'd9790256; ROM4[2955]<=26'd23533365;
ROM1[2956]<=26'd2164761; ROM2[2956]<=26'd11377107; ROM3[2956]<=26'd9784057; ROM4[2956]<=26'd23529670;
ROM1[2957]<=26'd2167322; ROM2[2957]<=26'd11372075; ROM3[2957]<=26'd9774180; ROM4[2957]<=26'd23522128;
ROM1[2958]<=26'd2166171; ROM2[2958]<=26'd11367507; ROM3[2958]<=26'd9768677; ROM4[2958]<=26'd23517018;
ROM1[2959]<=26'd2156681; ROM2[2959]<=26'd11366049; ROM3[2959]<=26'd9769100; ROM4[2959]<=26'd23516289;
ROM1[2960]<=26'd2145282; ROM2[2960]<=26'd11364267; ROM3[2960]<=26'd9771534; ROM4[2960]<=26'd23515502;
ROM1[2961]<=26'd2140211; ROM2[2961]<=26'd11367832; ROM3[2961]<=26'd9780058; ROM4[2961]<=26'd23520403;
ROM1[2962]<=26'd2126885; ROM2[2962]<=26'd11364896; ROM3[2962]<=26'd9778817; ROM4[2962]<=26'd23518320;
ROM1[2963]<=26'd2119754; ROM2[2963]<=26'd11362254; ROM3[2963]<=26'd9779214; ROM4[2963]<=26'd23516470;
ROM1[2964]<=26'd2119996; ROM2[2964]<=26'd11362626; ROM3[2964]<=26'd9780248; ROM4[2964]<=26'd23517866;
ROM1[2965]<=26'd2117159; ROM2[2965]<=26'd11351319; ROM3[2965]<=26'd9764376; ROM4[2965]<=26'd23506801;
ROM1[2966]<=26'd2122129; ROM2[2966]<=26'd11348770; ROM3[2966]<=26'd9754857; ROM4[2966]<=26'd23501287;
ROM1[2967]<=26'd2123245; ROM2[2967]<=26'd11354517; ROM3[2967]<=26'd9759292; ROM4[2967]<=26'd23506885;
ROM1[2968]<=26'd2112762; ROM2[2968]<=26'd11352289; ROM3[2968]<=26'd9761992; ROM4[2968]<=26'd23508050;
ROM1[2969]<=26'd2102459; ROM2[2969]<=26'd11351116; ROM3[2969]<=26'd9765251; ROM4[2969]<=26'd23508405;
ROM1[2970]<=26'd2097359; ROM2[2970]<=26'd11353179; ROM3[2970]<=26'd9771939; ROM4[2970]<=26'd23512107;
ROM1[2971]<=26'd2086800; ROM2[2971]<=26'd11349271; ROM3[2971]<=26'd9773365; ROM4[2971]<=26'd23510033;
ROM1[2972]<=26'd2082882; ROM2[2972]<=26'd11346238; ROM3[2972]<=26'd9770001; ROM4[2972]<=26'd23507208;
ROM1[2973]<=26'd2089896; ROM2[2973]<=26'd11348156; ROM3[2973]<=26'd9766441; ROM4[2973]<=26'd23506144;
ROM1[2974]<=26'd2097292; ROM2[2974]<=26'd11345458; ROM3[2974]<=26'd9760150; ROM4[2974]<=26'd23502106;
ROM1[2975]<=26'd2093132; ROM2[2975]<=26'd11339040; ROM3[2975]<=26'd9754105; ROM4[2975]<=26'd23498048;
ROM1[2976]<=26'd2081307; ROM2[2976]<=26'd11335562; ROM3[2976]<=26'd9754777; ROM4[2976]<=26'd23495346;
ROM1[2977]<=26'd2072713; ROM2[2977]<=26'd11335748; ROM3[2977]<=26'd9760805; ROM4[2977]<=26'd23497077;
ROM1[2978]<=26'd2071071; ROM2[2978]<=26'd11340324; ROM3[2978]<=26'd9770325; ROM4[2978]<=26'd23504948;
ROM1[2979]<=26'd2067544; ROM2[2979]<=26'd11345549; ROM3[2979]<=26'd9777819; ROM4[2979]<=26'd23508560;
ROM1[2980]<=26'd2056268; ROM2[2980]<=26'd11338691; ROM3[2980]<=26'd9769439; ROM4[2980]<=26'd23499271;
ROM1[2981]<=26'd2056895; ROM2[2981]<=26'd11335013; ROM3[2981]<=26'd9761238; ROM4[2981]<=26'd23494139;
ROM1[2982]<=26'd2067664; ROM2[2982]<=26'd11336284; ROM3[2982]<=26'd9755596; ROM4[2982]<=26'd23492021;
ROM1[2983]<=26'd2067713; ROM2[2983]<=26'd11331236; ROM3[2983]<=26'd9746106; ROM4[2983]<=26'd23486618;
ROM1[2984]<=26'd2062538; ROM2[2984]<=26'd11331378; ROM3[2984]<=26'd9748568; ROM4[2984]<=26'd23489071;
ROM1[2985]<=26'd2054003; ROM2[2985]<=26'd11332964; ROM3[2985]<=26'd9754333; ROM4[2985]<=26'd23490499;
ROM1[2986]<=26'd2045018; ROM2[2986]<=26'd11330049; ROM3[2986]<=26'd9755350; ROM4[2986]<=26'd23488868;
ROM1[2987]<=26'd2037750; ROM2[2987]<=26'd11328858; ROM3[2987]<=26'd9759411; ROM4[2987]<=26'd23490916;
ROM1[2988]<=26'd2034719; ROM2[2988]<=26'd11330947; ROM3[2988]<=26'd9763581; ROM4[2988]<=26'd23492885;
ROM1[2989]<=26'd2042300; ROM2[2989]<=26'd11334408; ROM3[2989]<=26'd9767105; ROM4[2989]<=26'd23496711;
ROM1[2990]<=26'd2053550; ROM2[2990]<=26'd11337125; ROM3[2990]<=26'd9765236; ROM4[2990]<=26'd23498373;
ROM1[2991]<=26'd2064459; ROM2[2991]<=26'd11339720; ROM3[2991]<=26'd9760811; ROM4[2991]<=26'd23497413;
ROM1[2992]<=26'd2068105; ROM2[2992]<=26'd11344105; ROM3[2992]<=26'd9767721; ROM4[2992]<=26'd23502746;
ROM1[2993]<=26'd2053113; ROM2[2993]<=26'd11337188; ROM3[2993]<=26'd9767015; ROM4[2993]<=26'd23499076;
ROM1[2994]<=26'd2039923; ROM2[2994]<=26'd11331423; ROM3[2994]<=26'd9765788; ROM4[2994]<=26'd23496177;
ROM1[2995]<=26'd2035107; ROM2[2995]<=26'd11329914; ROM3[2995]<=26'd9768543; ROM4[2995]<=26'd23496919;
ROM1[2996]<=26'd2023865; ROM2[2996]<=26'd11324036; ROM3[2996]<=26'd9764504; ROM4[2996]<=26'd23489417;
ROM1[2997]<=26'd2024026; ROM2[2997]<=26'd11325286; ROM3[2997]<=26'd9762858; ROM4[2997]<=26'd23488421;
ROM1[2998]<=26'd2037363; ROM2[2998]<=26'd11329727; ROM3[2998]<=26'd9763303; ROM4[2998]<=26'd23489531;
ROM1[2999]<=26'd2052563; ROM2[2999]<=26'd11335297; ROM3[2999]<=26'd9761457; ROM4[2999]<=26'd23491827;
ROM1[3000]<=26'd2053076; ROM2[3000]<=26'd11335404; ROM3[3000]<=26'd9758960; ROM4[3000]<=26'd23490533;
ROM1[3001]<=26'd2042282; ROM2[3001]<=26'd11329575; ROM3[3001]<=26'd9755365; ROM4[3001]<=26'd23485252;
ROM1[3002]<=26'd2032276; ROM2[3002]<=26'd11328002; ROM3[3002]<=26'd9755619; ROM4[3002]<=26'd23483934;
ROM1[3003]<=26'd2027026; ROM2[3003]<=26'd11328996; ROM3[3003]<=26'd9759032; ROM4[3003]<=26'd23484980;
ROM1[3004]<=26'd2025334; ROM2[3004]<=26'd11332392; ROM3[3004]<=26'd9764957; ROM4[3004]<=26'd23490150;
ROM1[3005]<=26'd2027586; ROM2[3005]<=26'd11336517; ROM3[3005]<=26'd9771744; ROM4[3005]<=26'd23493509;
ROM1[3006]<=26'd2027411; ROM2[3006]<=26'd11331248; ROM3[3006]<=26'd9764747; ROM4[3006]<=26'd23487879;
ROM1[3007]<=26'd2031077; ROM2[3007]<=26'd11324783; ROM3[3007]<=26'd9751523; ROM4[3007]<=26'd23479652;
ROM1[3008]<=26'd2029382; ROM2[3008]<=26'd11316451; ROM3[3008]<=26'd9740255; ROM4[3008]<=26'd23469853;
ROM1[3009]<=26'd2017281; ROM2[3009]<=26'd11310923; ROM3[3009]<=26'd9735306; ROM4[3009]<=26'd23463491;
ROM1[3010]<=26'd2008694; ROM2[3010]<=26'd11310391; ROM3[3010]<=26'd9735337; ROM4[3010]<=26'd23461243;
ROM1[3011]<=26'd2001336; ROM2[3011]<=26'd11307897; ROM3[3011]<=26'd9735104; ROM4[3011]<=26'd23457878;
ROM1[3012]<=26'd1992053; ROM2[3012]<=26'd11306775; ROM3[3012]<=26'd9735972; ROM4[3012]<=26'd23456616;
ROM1[3013]<=26'd1990442; ROM2[3013]<=26'd11307204; ROM3[3013]<=26'd9738700; ROM4[3013]<=26'd23458902;
ROM1[3014]<=26'd1998783; ROM2[3014]<=26'd11313649; ROM3[3014]<=26'd9741866; ROM4[3014]<=26'd23463368;
ROM1[3015]<=26'd2005446; ROM2[3015]<=26'd11312609; ROM3[3015]<=26'd9735036; ROM4[3015]<=26'd23459619;
ROM1[3016]<=26'd2009567; ROM2[3016]<=26'd11307214; ROM3[3016]<=26'd9727361; ROM4[3016]<=26'd23454683;
ROM1[3017]<=26'd2009552; ROM2[3017]<=26'd11310685; ROM3[3017]<=26'd9730989; ROM4[3017]<=26'd23458393;
ROM1[3018]<=26'd2003435; ROM2[3018]<=26'd11311488; ROM3[3018]<=26'd9737054; ROM4[3018]<=26'd23463411;
ROM1[3019]<=26'd2000072; ROM2[3019]<=26'd11312613; ROM3[3019]<=26'd9744723; ROM4[3019]<=26'd23468288;
ROM1[3020]<=26'd1996196; ROM2[3020]<=26'd11312131; ROM3[3020]<=26'd9747192; ROM4[3020]<=26'd23469145;
ROM1[3021]<=26'd1991492; ROM2[3021]<=26'd11312180; ROM3[3021]<=26'd9750190; ROM4[3021]<=26'd23469309;
ROM1[3022]<=26'd1997555; ROM2[3022]<=26'd11316887; ROM3[3022]<=26'd9756724; ROM4[3022]<=26'd23474530;
ROM1[3023]<=26'd2005036; ROM2[3023]<=26'd11318658; ROM3[3023]<=26'd9753652; ROM4[3023]<=26'd23474908;
ROM1[3024]<=26'd2018201; ROM2[3024]<=26'd11322249; ROM3[3024]<=26'd9750990; ROM4[3024]<=26'd23476712;
ROM1[3025]<=26'd2020227; ROM2[3025]<=26'd11321305; ROM3[3025]<=26'd9748010; ROM4[3025]<=26'd23476714;
ROM1[3026]<=26'd2007982; ROM2[3026]<=26'd11315072; ROM3[3026]<=26'd9744096; ROM4[3026]<=26'd23470421;
ROM1[3027]<=26'd1998199; ROM2[3027]<=26'd11313980; ROM3[3027]<=26'd9746108; ROM4[3027]<=26'd23468568;
ROM1[3028]<=26'd1994081; ROM2[3028]<=26'd11316296; ROM3[3028]<=26'd9748892; ROM4[3028]<=26'd23469656;
ROM1[3029]<=26'd1987293; ROM2[3029]<=26'd11314304; ROM3[3029]<=26'd9750113; ROM4[3029]<=26'd23467189;
ROM1[3030]<=26'd1981534; ROM2[3030]<=26'd11311238; ROM3[3030]<=26'd9746144; ROM4[3030]<=26'd23463373;
ROM1[3031]<=26'd1988815; ROM2[3031]<=26'd11311728; ROM3[3031]<=26'd9743846; ROM4[3031]<=26'd23462949;
ROM1[3032]<=26'd2003282; ROM2[3032]<=26'd11314860; ROM3[3032]<=26'd9742620; ROM4[3032]<=26'd23465139;
ROM1[3033]<=26'd2009189; ROM2[3033]<=26'd11315253; ROM3[3033]<=26'd9739106; ROM4[3033]<=26'd23466168;
ROM1[3034]<=26'd2007069; ROM2[3034]<=26'd11314390; ROM3[3034]<=26'd9743037; ROM4[3034]<=26'd23467295;
ROM1[3035]<=26'd2002999; ROM2[3035]<=26'd11315973; ROM3[3035]<=26'd9752065; ROM4[3035]<=26'd23471619;
ROM1[3036]<=26'd2001345; ROM2[3036]<=26'd11317676; ROM3[3036]<=26'd9759096; ROM4[3036]<=26'd23475329;
ROM1[3037]<=26'd1996780; ROM2[3037]<=26'd11316351; ROM3[3037]<=26'd9763729; ROM4[3037]<=26'd23475358;
ROM1[3038]<=26'd1995303; ROM2[3038]<=26'd11317060; ROM3[3038]<=26'd9766402; ROM4[3038]<=26'd23478453;
ROM1[3039]<=26'd2002293; ROM2[3039]<=26'd11319061; ROM3[3039]<=26'd9767899; ROM4[3039]<=26'd23482544;
ROM1[3040]<=26'd2014332; ROM2[3040]<=26'd11318805; ROM3[3040]<=26'd9764955; ROM4[3040]<=26'd23482781;
ROM1[3041]<=26'd2021430; ROM2[3041]<=26'd11317261; ROM3[3041]<=26'd9756583; ROM4[3041]<=26'd23478475;
ROM1[3042]<=26'd2014662; ROM2[3042]<=26'd11313100; ROM3[3042]<=26'd9752413; ROM4[3042]<=26'd23472976;
ROM1[3043]<=26'd2004271; ROM2[3043]<=26'd11309702; ROM3[3043]<=26'd9752273; ROM4[3043]<=26'd23470337;
ROM1[3044]<=26'd2000751; ROM2[3044]<=26'd11311318; ROM3[3044]<=26'd9757022; ROM4[3044]<=26'd23473150;
ROM1[3045]<=26'd2007224; ROM2[3045]<=26'd11322886; ROM3[3045]<=26'd9770188; ROM4[3045]<=26'd23486244;
ROM1[3046]<=26'd2010611; ROM2[3046]<=26'd11331736; ROM3[3046]<=26'd9780716; ROM4[3046]<=26'd23494350;
ROM1[3047]<=26'd2002427; ROM2[3047]<=26'd11322520; ROM3[3047]<=26'd9771599; ROM4[3047]<=26'd23484894;
ROM1[3048]<=26'd1997821; ROM2[3048]<=26'd11311683; ROM3[3048]<=26'd9755758; ROM4[3048]<=26'd23472312;
ROM1[3049]<=26'd2008875; ROM2[3049]<=26'd11312508; ROM3[3049]<=26'd9751728; ROM4[3049]<=26'd23472008;
ROM1[3050]<=26'd2007134; ROM2[3050]<=26'd11308859; ROM3[3050]<=26'd9750913; ROM4[3050]<=26'd23472131;
ROM1[3051]<=26'd2001490; ROM2[3051]<=26'd11310153; ROM3[3051]<=26'd9753793; ROM4[3051]<=26'd23475341;
ROM1[3052]<=26'd1998354; ROM2[3052]<=26'd11315569; ROM3[3052]<=26'd9760084; ROM4[3052]<=26'd23480096;
ROM1[3053]<=26'd1985881; ROM2[3053]<=26'd11308519; ROM3[3053]<=26'd9756849; ROM4[3053]<=26'd23476716;
ROM1[3054]<=26'd1974024; ROM2[3054]<=26'd11304430; ROM3[3054]<=26'd9754061; ROM4[3054]<=26'd23474067;
ROM1[3055]<=26'd1977020; ROM2[3055]<=26'd11310871; ROM3[3055]<=26'd9760669; ROM4[3055]<=26'd23478682;
ROM1[3056]<=26'd1987875; ROM2[3056]<=26'd11317257; ROM3[3056]<=26'd9764440; ROM4[3056]<=26'd23484501;
ROM1[3057]<=26'd1987344; ROM2[3057]<=26'd11306650; ROM3[3057]<=26'd9745885; ROM4[3057]<=26'd23471808;
ROM1[3058]<=26'd1985446; ROM2[3058]<=26'd11296985; ROM3[3058]<=26'd9731681; ROM4[3058]<=26'd23461018;
ROM1[3059]<=26'd1981955; ROM2[3059]<=26'd11295574; ROM3[3059]<=26'd9730802; ROM4[3059]<=26'd23459323;
ROM1[3060]<=26'd1972320; ROM2[3060]<=26'd11293031; ROM3[3060]<=26'd9731357; ROM4[3060]<=26'd23457728;
ROM1[3061]<=26'd1969389; ROM2[3061]<=26'd11295619; ROM3[3061]<=26'd9738048; ROM4[3061]<=26'd23460861;
ROM1[3062]<=26'd1972718; ROM2[3062]<=26'd11302194; ROM3[3062]<=26'd9746853; ROM4[3062]<=26'd23466563;
ROM1[3063]<=26'd1972392; ROM2[3063]<=26'd11303703; ROM3[3063]<=26'd9752148; ROM4[3063]<=26'd23469145;
ROM1[3064]<=26'd1970603; ROM2[3064]<=26'd11298437; ROM3[3064]<=26'd9745753; ROM4[3064]<=26'd23462731;
ROM1[3065]<=26'd1984230; ROM2[3065]<=26'd11300878; ROM3[3065]<=26'd9740857; ROM4[3065]<=26'd23461493;
ROM1[3066]<=26'd1999136; ROM2[3066]<=26'd11305121; ROM3[3066]<=26'd9740291; ROM4[3066]<=26'd23464312;
ROM1[3067]<=26'd1992915; ROM2[3067]<=26'd11299537; ROM3[3067]<=26'd9734791; ROM4[3067]<=26'd23457328;
ROM1[3068]<=26'd1985802; ROM2[3068]<=26'd11296679; ROM3[3068]<=26'd9737444; ROM4[3068]<=26'd23456523;
ROM1[3069]<=26'd1982852; ROM2[3069]<=26'd11296536; ROM3[3069]<=26'd9744810; ROM4[3069]<=26'd23459825;
ROM1[3070]<=26'd1974505; ROM2[3070]<=26'd11293884; ROM3[3070]<=26'd9745270; ROM4[3070]<=26'd23456472;
ROM1[3071]<=26'd1971285; ROM2[3071]<=26'd11294120; ROM3[3071]<=26'd9748463; ROM4[3071]<=26'd23458282;
ROM1[3072]<=26'd1975872; ROM2[3072]<=26'd11296780; ROM3[3072]<=26'd9750657; ROM4[3072]<=26'd23460813;
ROM1[3073]<=26'd1986405; ROM2[3073]<=26'd11299675; ROM3[3073]<=26'd9750453; ROM4[3073]<=26'd23462534;
ROM1[3074]<=26'd1996821; ROM2[3074]<=26'd11295977; ROM3[3074]<=26'd9747699; ROM4[3074]<=26'd23462511;
ROM1[3075]<=26'd1991454; ROM2[3075]<=26'd11286198; ROM3[3075]<=26'd9741932; ROM4[3075]<=26'd23455829;
ROM1[3076]<=26'd1986058; ROM2[3076]<=26'd11285469; ROM3[3076]<=26'd9746963; ROM4[3076]<=26'd23456919;
ROM1[3077]<=26'd1979824; ROM2[3077]<=26'd11284565; ROM3[3077]<=26'd9752238; ROM4[3077]<=26'd23457853;
ROM1[3078]<=26'd1971002; ROM2[3078]<=26'd11280871; ROM3[3078]<=26'd9752400; ROM4[3078]<=26'd23453580;
ROM1[3079]<=26'd1961232; ROM2[3079]<=26'd11278270; ROM3[3079]<=26'd9751810; ROM4[3079]<=26'd23449720;
ROM1[3080]<=26'd1955966; ROM2[3080]<=26'd11276156; ROM3[3080]<=26'd9748507; ROM4[3080]<=26'd23445338;
ROM1[3081]<=26'd1963029; ROM2[3081]<=26'd11279026; ROM3[3081]<=26'd9746407; ROM4[3081]<=26'd23445381;
ROM1[3082]<=26'd1982518; ROM2[3082]<=26'd11288730; ROM3[3082]<=26'd9745357; ROM4[3082]<=26'd23450930;
ROM1[3083]<=26'd1993327; ROM2[3083]<=26'd11295068; ROM3[3083]<=26'd9745302; ROM4[3083]<=26'd23455610;
ROM1[3084]<=26'd1976873; ROM2[3084]<=26'd11281496; ROM3[3084]<=26'd9735885; ROM4[3084]<=26'd23446241;
ROM1[3085]<=26'd1962582; ROM2[3085]<=26'd11272715; ROM3[3085]<=26'd9732275; ROM4[3085]<=26'd23440060;
ROM1[3086]<=26'd1960426; ROM2[3086]<=26'd11275525; ROM3[3086]<=26'd9738842; ROM4[3086]<=26'd23443933;
ROM1[3087]<=26'd1958270; ROM2[3087]<=26'd11279045; ROM3[3087]<=26'd9746697; ROM4[3087]<=26'd23451200;
ROM1[3088]<=26'd1964419; ROM2[3088]<=26'd11287508; ROM3[3088]<=26'd9757497; ROM4[3088]<=26'd23462662;
ROM1[3089]<=26'd1974655; ROM2[3089]<=26'd11293396; ROM3[3089]<=26'd9762682; ROM4[3089]<=26'd23469435;
ROM1[3090]<=26'd1983266; ROM2[3090]<=26'd11293529; ROM3[3090]<=26'd9758452; ROM4[3090]<=26'd23469790;
ROM1[3091]<=26'd1994471; ROM2[3091]<=26'd11295513; ROM3[3091]<=26'd9756366; ROM4[3091]<=26'd23473304;
ROM1[3092]<=26'd1998228; ROM2[3092]<=26'd11301496; ROM3[3092]<=26'd9760615; ROM4[3092]<=26'd23479613;
ROM1[3093]<=26'd1996467; ROM2[3093]<=26'd11306201; ROM3[3093]<=26'd9767943; ROM4[3093]<=26'd23486499;
ROM1[3094]<=26'd1989302; ROM2[3094]<=26'd11303227; ROM3[3094]<=26'd9771187; ROM4[3094]<=26'd23486657;
ROM1[3095]<=26'd1980417; ROM2[3095]<=26'd11299205; ROM3[3095]<=26'd9769410; ROM4[3095]<=26'd23482632;
ROM1[3096]<=26'd1977779; ROM2[3096]<=26'd11303052; ROM3[3096]<=26'd9772653; ROM4[3096]<=26'd23484701;
ROM1[3097]<=26'd1980179; ROM2[3097]<=26'd11305694; ROM3[3097]<=26'd9772802; ROM4[3097]<=26'd23485768;
ROM1[3098]<=26'd1992729; ROM2[3098]<=26'd11310631; ROM3[3098]<=26'd9768976; ROM4[3098]<=26'd23488027;
ROM1[3099]<=26'd2007205; ROM2[3099]<=26'd11314829; ROM3[3099]<=26'd9763165; ROM4[3099]<=26'd23487268;
ROM1[3100]<=26'd2006435; ROM2[3100]<=26'd11312171; ROM3[3100]<=26'd9759085; ROM4[3100]<=26'd23483481;
ROM1[3101]<=26'd1999019; ROM2[3101]<=26'd11312295; ROM3[3101]<=26'd9759682; ROM4[3101]<=26'd23482680;
ROM1[3102]<=26'd1988188; ROM2[3102]<=26'd11310104; ROM3[3102]<=26'd9759751; ROM4[3102]<=26'd23479489;
ROM1[3103]<=26'd1986477; ROM2[3103]<=26'd11313776; ROM3[3103]<=26'd9764104; ROM4[3103]<=26'd23481786;
ROM1[3104]<=26'd1986690; ROM2[3104]<=26'd11319253; ROM3[3104]<=26'd9768276; ROM4[3104]<=26'd23486077;
ROM1[3105]<=26'd1984340; ROM2[3105]<=26'd11319629; ROM3[3105]<=26'd9767567; ROM4[3105]<=26'd23483236;
ROM1[3106]<=26'd1988533; ROM2[3106]<=26'd11320226; ROM3[3106]<=26'd9761915; ROM4[3106]<=26'd23480530;
ROM1[3107]<=26'd1997755; ROM2[3107]<=26'd11317746; ROM3[3107]<=26'd9750769; ROM4[3107]<=26'd23476140;
ROM1[3108]<=26'd1998685; ROM2[3108]<=26'd11313346; ROM3[3108]<=26'd9742674; ROM4[3108]<=26'd23469022;
ROM1[3109]<=26'd1989025; ROM2[3109]<=26'd11308617; ROM3[3109]<=26'd9739556; ROM4[3109]<=26'd23465106;
ROM1[3110]<=26'd1981000; ROM2[3110]<=26'd11306721; ROM3[3110]<=26'd9742035; ROM4[3110]<=26'd23464099;
ROM1[3111]<=26'd1978463; ROM2[3111]<=26'd11308591; ROM3[3111]<=26'd9749230; ROM4[3111]<=26'd23466451;
ROM1[3112]<=26'd1972837; ROM2[3112]<=26'd11307240; ROM3[3112]<=26'd9752456; ROM4[3112]<=26'd23467389;
ROM1[3113]<=26'd1966750; ROM2[3113]<=26'd11303553; ROM3[3113]<=26'd9751083; ROM4[3113]<=26'd23464275;
ROM1[3114]<=26'd1969651; ROM2[3114]<=26'd11301941; ROM3[3114]<=26'd9748396; ROM4[3114]<=26'd23460957;
ROM1[3115]<=26'd1979846; ROM2[3115]<=26'd11301187; ROM3[3115]<=26'd9742974; ROM4[3115]<=26'd23458536;
ROM1[3116]<=26'd1993291; ROM2[3116]<=26'd11305645; ROM3[3116]<=26'd9741159; ROM4[3116]<=26'd23460077;
ROM1[3117]<=26'd1995905; ROM2[3117]<=26'd11309045; ROM3[3117]<=26'd9744516; ROM4[3117]<=26'd23462683;
ROM1[3118]<=26'd1984628; ROM2[3118]<=26'd11304201; ROM3[3118]<=26'd9742509; ROM4[3118]<=26'd23459286;
ROM1[3119]<=26'd1971522; ROM2[3119]<=26'd11297985; ROM3[3119]<=26'd9739469; ROM4[3119]<=26'd23454869;
ROM1[3120]<=26'd1972458; ROM2[3120]<=26'd11302792; ROM3[3120]<=26'd9747929; ROM4[3120]<=26'd23460574;
ROM1[3121]<=26'd1968541; ROM2[3121]<=26'd11302310; ROM3[3121]<=26'd9749808; ROM4[3121]<=26'd23461670;
ROM1[3122]<=26'd1963345; ROM2[3122]<=26'd11296533; ROM3[3122]<=26'd9744920; ROM4[3122]<=26'd23456217;
ROM1[3123]<=26'd1969696; ROM2[3123]<=26'd11295218; ROM3[3123]<=26'd9739443; ROM4[3123]<=26'd23453671;
ROM1[3124]<=26'd1982236; ROM2[3124]<=26'd11296270; ROM3[3124]<=26'd9734736; ROM4[3124]<=26'd23454569;
ROM1[3125]<=26'd1985287; ROM2[3125]<=26'd11296329; ROM3[3125]<=26'd9733707; ROM4[3125]<=26'd23455005;
ROM1[3126]<=26'd1981751; ROM2[3126]<=26'd11296552; ROM3[3126]<=26'd9738150; ROM4[3126]<=26'd23456512;
ROM1[3127]<=26'd1978241; ROM2[3127]<=26'd11299919; ROM3[3127]<=26'd9745707; ROM4[3127]<=26'd23461123;
ROM1[3128]<=26'd1970030; ROM2[3128]<=26'd11296832; ROM3[3128]<=26'd9745136; ROM4[3128]<=26'd23459333;
ROM1[3129]<=26'd1965618; ROM2[3129]<=26'd11295348; ROM3[3129]<=26'd9747620; ROM4[3129]<=26'd23459645;
ROM1[3130]<=26'd1970174; ROM2[3130]<=26'd11301854; ROM3[3130]<=26'd9752652; ROM4[3130]<=26'd23466744;
ROM1[3131]<=26'd1980618; ROM2[3131]<=26'd11306041; ROM3[3131]<=26'd9753447; ROM4[3131]<=26'd23470542;
ROM1[3132]<=26'd1993380; ROM2[3132]<=26'd11307124; ROM3[3132]<=26'd9748846; ROM4[3132]<=26'd23470689;
ROM1[3133]<=26'd2006160; ROM2[3133]<=26'd11315421; ROM3[3133]<=26'd9754250; ROM4[3133]<=26'd23478242;
ROM1[3134]<=26'd2006865; ROM2[3134]<=26'd11319437; ROM3[3134]<=26'd9761862; ROM4[3134]<=26'd23485293;
ROM1[3135]<=26'd1999219; ROM2[3135]<=26'd11317848; ROM3[3135]<=26'd9764742; ROM4[3135]<=26'd23487226;
ROM1[3136]<=26'd1992190; ROM2[3136]<=26'd11312948; ROM3[3136]<=26'd9765155; ROM4[3136]<=26'd23485042;
ROM1[3137]<=26'd1982870; ROM2[3137]<=26'd11308229; ROM3[3137]<=26'd9764564; ROM4[3137]<=26'd23482922;
ROM1[3138]<=26'd1978000; ROM2[3138]<=26'd11308075; ROM3[3138]<=26'd9765633; ROM4[3138]<=26'd23483141;
ROM1[3139]<=26'd1983315; ROM2[3139]<=26'd11310431; ROM3[3139]<=26'd9766117; ROM4[3139]<=26'd23485410;
ROM1[3140]<=26'd2001174; ROM2[3140]<=26'd11319518; ROM3[3140]<=26'd9769311; ROM4[3140]<=26'd23492311;
ROM1[3141]<=26'd2011804; ROM2[3141]<=26'd11319566; ROM3[3141]<=26'd9762179; ROM4[3141]<=26'd23491360;
ROM1[3142]<=26'd2002645; ROM2[3142]<=26'd11308202; ROM3[3142]<=26'd9752067; ROM4[3142]<=26'd23482163;
ROM1[3143]<=26'd1993641; ROM2[3143]<=26'd11304972; ROM3[3143]<=26'd9754259; ROM4[3143]<=26'd23480136;
ROM1[3144]<=26'd1983724; ROM2[3144]<=26'd11302006; ROM3[3144]<=26'd9755049; ROM4[3144]<=26'd23478450;
ROM1[3145]<=26'd1973704; ROM2[3145]<=26'd11297537; ROM3[3145]<=26'd9754632; ROM4[3145]<=26'd23475003;
ROM1[3146]<=26'd1970961; ROM2[3146]<=26'd11299667; ROM3[3146]<=26'd9758720; ROM4[3146]<=26'd23475561;
ROM1[3147]<=26'd1974489; ROM2[3147]<=26'd11300549; ROM3[3147]<=26'd9760654; ROM4[3147]<=26'd23475692;
ROM1[3148]<=26'd1981600; ROM2[3148]<=26'd11299963; ROM3[3148]<=26'd9756365; ROM4[3148]<=26'd23472687;
ROM1[3149]<=26'd1992396; ROM2[3149]<=26'd11301460; ROM3[3149]<=26'd9750554; ROM4[3149]<=26'd23471064;
ROM1[3150]<=26'd1992298; ROM2[3150]<=26'd11299716; ROM3[3150]<=26'd9746934; ROM4[3150]<=26'd23468774;
ROM1[3151]<=26'd1985355; ROM2[3151]<=26'd11302175; ROM3[3151]<=26'd9747449; ROM4[3151]<=26'd23467233;
ROM1[3152]<=26'd1977086; ROM2[3152]<=26'd11301292; ROM3[3152]<=26'd9750344; ROM4[3152]<=26'd23465130;
ROM1[3153]<=26'd1962600; ROM2[3153]<=26'd11291536; ROM3[3153]<=26'd9743569; ROM4[3153]<=26'd23454265;
ROM1[3154]<=26'd1956089; ROM2[3154]<=26'd11291663; ROM3[3154]<=26'd9742293; ROM4[3154]<=26'd23452279;
ROM1[3155]<=26'd1956786; ROM2[3155]<=26'd11293031; ROM3[3155]<=26'd9742601; ROM4[3155]<=26'd23453105;
ROM1[3156]<=26'd1960369; ROM2[3156]<=26'd11293120; ROM3[3156]<=26'd9735087; ROM4[3156]<=26'd23449709;
ROM1[3157]<=26'd1978617; ROM2[3157]<=26'd11302680; ROM3[3157]<=26'd9732832; ROM4[3157]<=26'd23454216;
ROM1[3158]<=26'd1994086; ROM2[3158]<=26'd11313131; ROM3[3158]<=26'd9737101; ROM4[3158]<=26'd23461512;
ROM1[3159]<=26'd1990005; ROM2[3159]<=26'd11316068; ROM3[3159]<=26'd9740160; ROM4[3159]<=26'd23463374;
ROM1[3160]<=26'd1973961; ROM2[3160]<=26'd11307844; ROM3[3160]<=26'd9736726; ROM4[3160]<=26'd23456584;
ROM1[3161]<=26'd1967551; ROM2[3161]<=26'd11306333; ROM3[3161]<=26'd9739723; ROM4[3161]<=26'd23457176;
ROM1[3162]<=26'd1962207; ROM2[3162]<=26'd11307778; ROM3[3162]<=26'd9743915; ROM4[3162]<=26'd23459019;
ROM1[3163]<=26'd1961144; ROM2[3163]<=26'd11307438; ROM3[3163]<=26'd9745170; ROM4[3163]<=26'd23459467;
ROM1[3164]<=26'd1972642; ROM2[3164]<=26'd11312578; ROM3[3164]<=26'd9747307; ROM4[3164]<=26'd23463414;
ROM1[3165]<=26'd1988211; ROM2[3165]<=26'd11318422; ROM3[3165]<=26'd9746041; ROM4[3165]<=26'd23466157;
ROM1[3166]<=26'd2000486; ROM2[3166]<=26'd11322085; ROM3[3166]<=26'd9743449; ROM4[3166]<=26'd23468200;
ROM1[3167]<=26'd1999529; ROM2[3167]<=26'd11322049; ROM3[3167]<=26'd9744108; ROM4[3167]<=26'd23469152;
ROM1[3168]<=26'd1993383; ROM2[3168]<=26'd11321922; ROM3[3168]<=26'd9747387; ROM4[3168]<=26'd23468656;
ROM1[3169]<=26'd1985059; ROM2[3169]<=26'd11317829; ROM3[3169]<=26'd9748704; ROM4[3169]<=26'd23465660;
ROM1[3170]<=26'd1977935; ROM2[3170]<=26'd11314192; ROM3[3170]<=26'd9748883; ROM4[3170]<=26'd23463421;
ROM1[3171]<=26'd1972466; ROM2[3171]<=26'd11311324; ROM3[3171]<=26'd9750462; ROM4[3171]<=26'd23461314;
ROM1[3172]<=26'd1975819; ROM2[3172]<=26'd11312883; ROM3[3172]<=26'd9751049; ROM4[3172]<=26'd23464075;
ROM1[3173]<=26'd1992138; ROM2[3173]<=26'd11320794; ROM3[3173]<=26'd9753944; ROM4[3173]<=26'd23472358;
ROM1[3174]<=26'd2004875; ROM2[3174]<=26'd11320588; ROM3[3174]<=26'd9748919; ROM4[3174]<=26'd23472539;
ROM1[3175]<=26'd1999453; ROM2[3175]<=26'd11312748; ROM3[3175]<=26'd9740807; ROM4[3175]<=26'd23466357;
ROM1[3176]<=26'd1994020; ROM2[3176]<=26'd11311174; ROM3[3176]<=26'd9744877; ROM4[3176]<=26'd23467346;
ROM1[3177]<=26'd1989085; ROM2[3177]<=26'd11311496; ROM3[3177]<=26'd9750223; ROM4[3177]<=26'd23468791;
ROM1[3178]<=26'd1980861; ROM2[3178]<=26'd11306843; ROM3[3178]<=26'd9751115; ROM4[3178]<=26'd23468057;
ROM1[3179]<=26'd1972938; ROM2[3179]<=26'd11304758; ROM3[3179]<=26'd9753539; ROM4[3179]<=26'd23467072;
ROM1[3180]<=26'd1969141; ROM2[3180]<=26'd11302490; ROM3[3180]<=26'd9751871; ROM4[3180]<=26'd23464913;
ROM1[3181]<=26'd1972893; ROM2[3181]<=26'd11299738; ROM3[3181]<=26'd9747259; ROM4[3181]<=26'd23462336;
ROM1[3182]<=26'd1985039; ROM2[3182]<=26'd11298541; ROM3[3182]<=26'd9742650; ROM4[3182]<=26'd23460051;
ROM1[3183]<=26'd1995313; ROM2[3183]<=26'd11301253; ROM3[3183]<=26'd9741819; ROM4[3183]<=26'd23462803;
ROM1[3184]<=26'd1991467; ROM2[3184]<=26'd11301620; ROM3[3184]<=26'd9744825; ROM4[3184]<=26'd23464720;
ROM1[3185]<=26'd1980153; ROM2[3185]<=26'd11296905; ROM3[3185]<=26'd9744654; ROM4[3185]<=26'd23460832;
ROM1[3186]<=26'd1976464; ROM2[3186]<=26'd11301879; ROM3[3186]<=26'd9747871; ROM4[3186]<=26'd23461997;
ROM1[3187]<=26'd1972718; ROM2[3187]<=26'd11302484; ROM3[3187]<=26'd9750996; ROM4[3187]<=26'd23462330;
ROM1[3188]<=26'd1973446; ROM2[3188]<=26'd11304603; ROM3[3188]<=26'd9756238; ROM4[3188]<=26'd23465603;
ROM1[3189]<=26'd1981165; ROM2[3189]<=26'd11309674; ROM3[3189]<=26'd9759293; ROM4[3189]<=26'd23471328;
ROM1[3190]<=26'd1984238; ROM2[3190]<=26'd11302238; ROM3[3190]<=26'd9748494; ROM4[3190]<=26'd23463689;
ROM1[3191]<=26'd1988638; ROM2[3191]<=26'd11298719; ROM3[3191]<=26'd9739122; ROM4[3191]<=26'd23458907;
ROM1[3192]<=26'd1987245; ROM2[3192]<=26'd11299922; ROM3[3192]<=26'd9738626; ROM4[3192]<=26'd23459850;
ROM1[3193]<=26'd1980169; ROM2[3193]<=26'd11300802; ROM3[3193]<=26'd9740280; ROM4[3193]<=26'd23457872;
ROM1[3194]<=26'd1980886; ROM2[3194]<=26'd11306664; ROM3[3194]<=26'd9749326; ROM4[3194]<=26'd23464835;
ROM1[3195]<=26'd1977140; ROM2[3195]<=26'd11307781; ROM3[3195]<=26'd9754459; ROM4[3195]<=26'd23467400;
ROM1[3196]<=26'd1965920; ROM2[3196]<=26'd11302638; ROM3[3196]<=26'd9749665; ROM4[3196]<=26'd23461818;
ROM1[3197]<=26'd1964791; ROM2[3197]<=26'd11299380; ROM3[3197]<=26'd9744706; ROM4[3197]<=26'd23457790;
ROM1[3198]<=26'd1980208; ROM2[3198]<=26'd11305352; ROM3[3198]<=26'd9746226; ROM4[3198]<=26'd23459496;
ROM1[3199]<=26'd2004351; ROM2[3199]<=26'd11318604; ROM3[3199]<=26'd9749913; ROM4[3199]<=26'd23469833;
ROM1[3200]<=26'd2002126; ROM2[3200]<=26'd11315367; ROM3[3200]<=26'd9742964; ROM4[3200]<=26'd23466343;
ROM1[3201]<=26'd1985398; ROM2[3201]<=26'd11304639; ROM3[3201]<=26'd9735502; ROM4[3201]<=26'd23458270;
ROM1[3202]<=26'd1976670; ROM2[3202]<=26'd11306004; ROM3[3202]<=26'd9740196; ROM4[3202]<=26'd23459888;
ROM1[3203]<=26'd1972858; ROM2[3203]<=26'd11306529; ROM3[3203]<=26'd9742422; ROM4[3203]<=26'd23460721;
ROM1[3204]<=26'd1974114; ROM2[3204]<=26'd11312863; ROM3[3204]<=26'd9748905; ROM4[3204]<=26'd23466023;
ROM1[3205]<=26'd1990762; ROM2[3205]<=26'd11328044; ROM3[3205]<=26'd9764506; ROM4[3205]<=26'd23481500;
ROM1[3206]<=26'd1998761; ROM2[3206]<=26'd11327120; ROM3[3206]<=26'd9761626; ROM4[3206]<=26'd23481435;
ROM1[3207]<=26'd1999489; ROM2[3207]<=26'd11318371; ROM3[3207]<=26'd9746169; ROM4[3207]<=26'd23470627;
ROM1[3208]<=26'd2002398; ROM2[3208]<=26'd11313464; ROM3[3208]<=26'd9740281; ROM4[3208]<=26'd23466672;
ROM1[3209]<=26'd1992799; ROM2[3209]<=26'd11308311; ROM3[3209]<=26'd9738135; ROM4[3209]<=26'd23461586;
ROM1[3210]<=26'd1983820; ROM2[3210]<=26'd11305674; ROM3[3210]<=26'd9739411; ROM4[3210]<=26'd23459992;
ROM1[3211]<=26'd1980538; ROM2[3211]<=26'd11306727; ROM3[3211]<=26'd9744835; ROM4[3211]<=26'd23461742;
ROM1[3212]<=26'd1978215; ROM2[3212]<=26'd11309220; ROM3[3212]<=26'd9753099; ROM4[3212]<=26'd23464386;
ROM1[3213]<=26'd1973281; ROM2[3213]<=26'd11308094; ROM3[3213]<=26'd9754876; ROM4[3213]<=26'd23463128;
ROM1[3214]<=26'd1976147; ROM2[3214]<=26'd11311010; ROM3[3214]<=26'd9752830; ROM4[3214]<=26'd23464839;
ROM1[3215]<=26'd1996123; ROM2[3215]<=26'd11320069; ROM3[3215]<=26'd9755983; ROM4[3215]<=26'd23472878;
ROM1[3216]<=26'd2004568; ROM2[3216]<=26'd11316607; ROM3[3216]<=26'd9748136; ROM4[3216]<=26'd23470043;
ROM1[3217]<=26'd1993169; ROM2[3217]<=26'd11306249; ROM3[3217]<=26'd9737330; ROM4[3217]<=26'd23461413;
ROM1[3218]<=26'd1985707; ROM2[3218]<=26'd11302670; ROM3[3218]<=26'd9737800; ROM4[3218]<=26'd23459445;
ROM1[3219]<=26'd1977794; ROM2[3219]<=26'd11299356; ROM3[3219]<=26'd9739081; ROM4[3219]<=26'd23457232;
ROM1[3220]<=26'd1973073; ROM2[3220]<=26'd11302445; ROM3[3220]<=26'd9742965; ROM4[3220]<=26'd23459578;
ROM1[3221]<=26'd1971297; ROM2[3221]<=26'd11306629; ROM3[3221]<=26'd9748395; ROM4[3221]<=26'd23462760;
ROM1[3222]<=26'd1970579; ROM2[3222]<=26'd11305118; ROM3[3222]<=26'd9746307; ROM4[3222]<=26'd23461022;
ROM1[3223]<=26'd1976449; ROM2[3223]<=26'd11304455; ROM3[3223]<=26'd9740358; ROM4[3223]<=26'd23458853;
ROM1[3224]<=26'd1987457; ROM2[3224]<=26'd11305039; ROM3[3224]<=26'd9736025; ROM4[3224]<=26'd23457377;
ROM1[3225]<=26'd1994753; ROM2[3225]<=26'd11310657; ROM3[3225]<=26'd9739682; ROM4[3225]<=26'd23463168;
ROM1[3226]<=26'd1990830; ROM2[3226]<=26'd11312911; ROM3[3226]<=26'd9743904; ROM4[3226]<=26'd23464738;
ROM1[3227]<=26'd1983453; ROM2[3227]<=26'd11313579; ROM3[3227]<=26'd9748156; ROM4[3227]<=26'd23465232;
ROM1[3228]<=26'd1986233; ROM2[3228]<=26'd11321192; ROM3[3228]<=26'd9757494; ROM4[3228]<=26'd23473800;
ROM1[3229]<=26'd1984736; ROM2[3229]<=26'd11324065; ROM3[3229]<=26'd9764406; ROM4[3229]<=26'd23476507;
ROM1[3230]<=26'd1974833; ROM2[3230]<=26'd11316289; ROM3[3230]<=26'd9756365; ROM4[3230]<=26'd23466464;
ROM1[3231]<=26'd1975343; ROM2[3231]<=26'd11311762; ROM3[3231]<=26'd9747559; ROM4[3231]<=26'd23459914;
ROM1[3232]<=26'd1987025; ROM2[3232]<=26'd11312518; ROM3[3232]<=26'd9740959; ROM4[3232]<=26'd23459112;
ROM1[3233]<=26'd1992672; ROM2[3233]<=26'd11314072; ROM3[3233]<=26'd9735867; ROM4[3233]<=26'd23458658;
ROM1[3234]<=26'd1995502; ROM2[3234]<=26'd11320267; ROM3[3234]<=26'd9741928; ROM4[3234]<=26'd23465784;
ROM1[3235]<=26'd1995569; ROM2[3235]<=26'd11324884; ROM3[3235]<=26'd9749497; ROM4[3235]<=26'd23472787;
ROM1[3236]<=26'd1990291; ROM2[3236]<=26'd11324649; ROM3[3236]<=26'd9752592; ROM4[3236]<=26'd23473528;
ROM1[3237]<=26'd1986910; ROM2[3237]<=26'd11326482; ROM3[3237]<=26'd9755729; ROM4[3237]<=26'd23475813;
ROM1[3238]<=26'd1988621; ROM2[3238]<=26'd11329805; ROM3[3238]<=26'd9761783; ROM4[3238]<=26'd23479395;
ROM1[3239]<=26'd1983324; ROM2[3239]<=26'd11321315; ROM3[3239]<=26'd9751998; ROM4[3239]<=26'd23469138;
ROM1[3240]<=26'd1984953; ROM2[3240]<=26'd11313132; ROM3[3240]<=26'd9737261; ROM4[3240]<=26'd23458986;
ROM1[3241]<=26'd1994048; ROM2[3241]<=26'd11312850; ROM3[3241]<=26'd9731816; ROM4[3241]<=26'd23457470;
ROM1[3242]<=26'd1991003; ROM2[3242]<=26'd11311688; ROM3[3242]<=26'd9731358; ROM4[3242]<=26'd23457840;
ROM1[3243]<=26'd1987550; ROM2[3243]<=26'd11314249; ROM3[3243]<=26'd9739420; ROM4[3243]<=26'd23464272;
ROM1[3244]<=26'd1986163; ROM2[3244]<=26'd11316743; ROM3[3244]<=26'd9747816; ROM4[3244]<=26'd23468759;
ROM1[3245]<=26'd1979624; ROM2[3245]<=26'd11312614; ROM3[3245]<=26'd9750166; ROM4[3245]<=26'd23466721;
ROM1[3246]<=26'd1973573; ROM2[3246]<=26'd11309613; ROM3[3246]<=26'd9751003; ROM4[3246]<=26'd23466528;
ROM1[3247]<=26'd1976166; ROM2[3247]<=26'd11310600; ROM3[3247]<=26'd9752413; ROM4[3247]<=26'd23468398;
ROM1[3248]<=26'd1986462; ROM2[3248]<=26'd11313399; ROM3[3248]<=26'd9749994; ROM4[3248]<=26'd23469595;
ROM1[3249]<=26'd1998276; ROM2[3249]<=26'd11313617; ROM3[3249]<=26'd9741695; ROM4[3249]<=26'd23467649;
ROM1[3250]<=26'd2001485; ROM2[3250]<=26'd11314654; ROM3[3250]<=26'd9741135; ROM4[3250]<=26'd23468965;
ROM1[3251]<=26'd1998918; ROM2[3251]<=26'd11318460; ROM3[3251]<=26'd9746968; ROM4[3251]<=26'd23473906;
ROM1[3252]<=26'd1988823; ROM2[3252]<=26'd11317572; ROM3[3252]<=26'd9749560; ROM4[3252]<=26'd23473051;
ROM1[3253]<=26'd1984704; ROM2[3253]<=26'd11318547; ROM3[3253]<=26'd9753453; ROM4[3253]<=26'd23475309;
ROM1[3254]<=26'd1973627; ROM2[3254]<=26'd11312557; ROM3[3254]<=26'd9749952; ROM4[3254]<=26'd23471149;
ROM1[3255]<=26'd1967918; ROM2[3255]<=26'd11306545; ROM3[3255]<=26'd9743812; ROM4[3255]<=26'd23464455;
ROM1[3256]<=26'd1979499; ROM2[3256]<=26'd11310395; ROM3[3256]<=26'd9743000; ROM4[3256]<=26'd23466451;
ROM1[3257]<=26'd1989611; ROM2[3257]<=26'd11309054; ROM3[3257]<=26'd9736417; ROM4[3257]<=26'd23463718;
ROM1[3258]<=26'd1999085; ROM2[3258]<=26'd11313231; ROM3[3258]<=26'd9735103; ROM4[3258]<=26'd23465443;
ROM1[3259]<=26'd1994739; ROM2[3259]<=26'd11312702; ROM3[3259]<=26'd9734642; ROM4[3259]<=26'd23463712;
ROM1[3260]<=26'd1982041; ROM2[3260]<=26'd11304903; ROM3[3260]<=26'd9732405; ROM4[3260]<=26'd23457606;
ROM1[3261]<=26'd1981197; ROM2[3261]<=26'd11311740; ROM3[3261]<=26'd9741705; ROM4[3261]<=26'd23464856;
ROM1[3262]<=26'd1972938; ROM2[3262]<=26'd11309778; ROM3[3262]<=26'd9742755; ROM4[3262]<=26'd23464622;
ROM1[3263]<=26'd1962568; ROM2[3263]<=26'd11299262; ROM3[3263]<=26'd9735669; ROM4[3263]<=26'd23455613;
ROM1[3264]<=26'd1970498; ROM2[3264]<=26'd11303188; ROM3[3264]<=26'd9736608; ROM4[3264]<=26'd23458581;
ROM1[3265]<=26'd1983551; ROM2[3265]<=26'd11305476; ROM3[3265]<=26'd9732595; ROM4[3265]<=26'd23458777;
ROM1[3266]<=26'd1995331; ROM2[3266]<=26'd11306657; ROM3[3266]<=26'd9730680; ROM4[3266]<=26'd23459480;
ROM1[3267]<=26'd1998373; ROM2[3267]<=26'd11315094; ROM3[3267]<=26'd9737343; ROM4[3267]<=26'd23467413;
ROM1[3268]<=26'd1991231; ROM2[3268]<=26'd11315327; ROM3[3268]<=26'd9739470; ROM4[3268]<=26'd23467834;
ROM1[3269]<=26'd1981799; ROM2[3269]<=26'd11310114; ROM3[3269]<=26'd9739204; ROM4[3269]<=26'd23465719;
ROM1[3270]<=26'd1977013; ROM2[3270]<=26'd11311749; ROM3[3270]<=26'd9741717; ROM4[3270]<=26'd23467344;
ROM1[3271]<=26'd1975763; ROM2[3271]<=26'd11314763; ROM3[3271]<=26'd9747914; ROM4[3271]<=26'd23469887;
ROM1[3272]<=26'd1979840; ROM2[3272]<=26'd11317098; ROM3[3272]<=26'd9751402; ROM4[3272]<=26'd23474309;
ROM1[3273]<=26'd1990904; ROM2[3273]<=26'd11319541; ROM3[3273]<=26'd9748343; ROM4[3273]<=26'd23476276;
ROM1[3274]<=26'd2004957; ROM2[3274]<=26'd11320929; ROM3[3274]<=26'd9744248; ROM4[3274]<=26'd23475803;
ROM1[3275]<=26'd2006547; ROM2[3275]<=26'd11321832; ROM3[3275]<=26'd9742954; ROM4[3275]<=26'd23476395;
ROM1[3276]<=26'd2002177; ROM2[3276]<=26'd11324162; ROM3[3276]<=26'd9746996; ROM4[3276]<=26'd23479086;
ROM1[3277]<=26'd1999112; ROM2[3277]<=26'd11327304; ROM3[3277]<=26'd9755608; ROM4[3277]<=26'd23483896;
ROM1[3278]<=26'd1992718; ROM2[3278]<=26'd11326951; ROM3[3278]<=26'd9759223; ROM4[3278]<=26'd23484191;
ROM1[3279]<=26'd1984155; ROM2[3279]<=26'd11322214; ROM3[3279]<=26'd9757297; ROM4[3279]<=26'd23479959;
ROM1[3280]<=26'd1982217; ROM2[3280]<=26'd11319557; ROM3[3280]<=26'd9755847; ROM4[3280]<=26'd23477173;
ROM1[3281]<=26'd1984091; ROM2[3281]<=26'd11316647; ROM3[3281]<=26'd9749906; ROM4[3281]<=26'd23472385;
ROM1[3282]<=26'd1995003; ROM2[3282]<=26'd11316487; ROM3[3282]<=26'd9744228; ROM4[3282]<=26'd23470573;
ROM1[3283]<=26'd2004781; ROM2[3283]<=26'd11317965; ROM3[3283]<=26'd9744433; ROM4[3283]<=26'd23473968;
ROM1[3284]<=26'd2000228; ROM2[3284]<=26'd11317970; ROM3[3284]<=26'd9746353; ROM4[3284]<=26'd23476096;
ROM1[3285]<=26'd1995074; ROM2[3285]<=26'd11319212; ROM3[3285]<=26'd9751870; ROM4[3285]<=26'd23479402;
ROM1[3286]<=26'd1993262; ROM2[3286]<=26'd11320942; ROM3[3286]<=26'd9757753; ROM4[3286]<=26'd23482915;
ROM1[3287]<=26'd1987473; ROM2[3287]<=26'd11321689; ROM3[3287]<=26'd9761951; ROM4[3287]<=26'd23482912;
ROM1[3288]<=26'd1979328; ROM2[3288]<=26'd11316852; ROM3[3288]<=26'd9761408; ROM4[3288]<=26'd23479952;
ROM1[3289]<=26'd1978846; ROM2[3289]<=26'd11313193; ROM3[3289]<=26'd9758094; ROM4[3289]<=26'd23475828;
ROM1[3290]<=26'd1991695; ROM2[3290]<=26'd11314918; ROM3[3290]<=26'd9753830; ROM4[3290]<=26'd23475506;
ROM1[3291]<=26'd2004567; ROM2[3291]<=26'd11318033; ROM3[3291]<=26'd9752296; ROM4[3291]<=26'd23479828;
ROM1[3292]<=26'd2001333; ROM2[3292]<=26'd11317821; ROM3[3292]<=26'd9753609; ROM4[3292]<=26'd23478749;
ROM1[3293]<=26'd1993736; ROM2[3293]<=26'd11316815; ROM3[3293]<=26'd9753473; ROM4[3293]<=26'd23476064;
ROM1[3294]<=26'd1987183; ROM2[3294]<=26'd11315816; ROM3[3294]<=26'd9755051; ROM4[3294]<=26'd23474844;
ROM1[3295]<=26'd1986281; ROM2[3295]<=26'd11322078; ROM3[3295]<=26'd9762502; ROM4[3295]<=26'd23477911;
ROM1[3296]<=26'd1983532; ROM2[3296]<=26'd11322542; ROM3[3296]<=26'd9761853; ROM4[3296]<=26'd23477166;
ROM1[3297]<=26'd1979268; ROM2[3297]<=26'd11315642; ROM3[3297]<=26'd9752380; ROM4[3297]<=26'd23469781;
ROM1[3298]<=26'd1990328; ROM2[3298]<=26'd11320812; ROM3[3298]<=26'd9750961; ROM4[3298]<=26'd23473003;
ROM1[3299]<=26'd2003769; ROM2[3299]<=26'd11324116; ROM3[3299]<=26'd9745435; ROM4[3299]<=26'd23474337;
ROM1[3300]<=26'd2004805; ROM2[3300]<=26'd11323183; ROM3[3300]<=26'd9743540; ROM4[3300]<=26'd23473056;
ROM1[3301]<=26'd1999427; ROM2[3301]<=26'd11325014; ROM3[3301]<=26'd9747371; ROM4[3301]<=26'd23474636;
ROM1[3302]<=26'd1990085; ROM2[3302]<=26'd11322295; ROM3[3302]<=26'd9748278; ROM4[3302]<=26'd23471811;
ROM1[3303]<=26'd1983082; ROM2[3303]<=26'd11316839; ROM3[3303]<=26'd9747175; ROM4[3303]<=26'd23468510;
ROM1[3304]<=26'd1979702; ROM2[3304]<=26'd11315934; ROM3[3304]<=26'd9749579; ROM4[3304]<=26'd23468264;
ROM1[3305]<=26'd1983915; ROM2[3305]<=26'd11318783; ROM3[3305]<=26'd9756052; ROM4[3305]<=26'd23472794;
ROM1[3306]<=26'd1992892; ROM2[3306]<=26'd11320441; ROM3[3306]<=26'd9755819; ROM4[3306]<=26'd23474292;
ROM1[3307]<=26'd2006341; ROM2[3307]<=26'd11320931; ROM3[3307]<=26'd9749975; ROM4[3307]<=26'd23472981;
ROM1[3308]<=26'd2009697; ROM2[3308]<=26'd11318280; ROM3[3308]<=26'd9745613; ROM4[3308]<=26'd23471259;
ROM1[3309]<=26'd2003353; ROM2[3309]<=26'd11315732; ROM3[3309]<=26'd9747107; ROM4[3309]<=26'd23470810;
ROM1[3310]<=26'd1999604; ROM2[3310]<=26'd11316697; ROM3[3310]<=26'd9753931; ROM4[3310]<=26'd23474606;
ROM1[3311]<=26'd1992046; ROM2[3311]<=26'd11313703; ROM3[3311]<=26'd9756822; ROM4[3311]<=26'd23474695;
ROM1[3312]<=26'd1984162; ROM2[3312]<=26'd11311467; ROM3[3312]<=26'd9756323; ROM4[3312]<=26'd23471730;
ROM1[3313]<=26'd1982476; ROM2[3313]<=26'd11314056; ROM3[3313]<=26'd9758817; ROM4[3313]<=26'd23471853;
ROM1[3314]<=26'd1986426; ROM2[3314]<=26'd11316211; ROM3[3314]<=26'd9757783; ROM4[3314]<=26'd23471161;
ROM1[3315]<=26'd1996516; ROM2[3315]<=26'd11316701; ROM3[3315]<=26'd9753326; ROM4[3315]<=26'd23470965;
ROM1[3316]<=26'd2003900; ROM2[3316]<=26'd11316025; ROM3[3316]<=26'd9749036; ROM4[3316]<=26'd23471072;
ROM1[3317]<=26'd2000930; ROM2[3317]<=26'd11314297; ROM3[3317]<=26'd9748967; ROM4[3317]<=26'd23470107;
ROM1[3318]<=26'd1990649; ROM2[3318]<=26'd11309847; ROM3[3318]<=26'd9749898; ROM4[3318]<=26'd23466266;
ROM1[3319]<=26'd1985171; ROM2[3319]<=26'd11308255; ROM3[3319]<=26'd9752075; ROM4[3319]<=26'd23463888;
ROM1[3320]<=26'd1987162; ROM2[3320]<=26'd11313937; ROM3[3320]<=26'd9759000; ROM4[3320]<=26'd23469294;
ROM1[3321]<=26'd1987922; ROM2[3321]<=26'd11318381; ROM3[3321]<=26'd9764440; ROM4[3321]<=26'd23474196;
ROM1[3322]<=26'd1991915; ROM2[3322]<=26'd11319931; ROM3[3322]<=26'd9765154; ROM4[3322]<=26'd23477767;
ROM1[3323]<=26'd1994349; ROM2[3323]<=26'd11316160; ROM3[3323]<=26'd9754911; ROM4[3323]<=26'd23472136;
ROM1[3324]<=26'd2003941; ROM2[3324]<=26'd11315914; ROM3[3324]<=26'd9745433; ROM4[3324]<=26'd23467414;
ROM1[3325]<=26'd2009857; ROM2[3325]<=26'd11318936; ROM3[3325]<=26'd9745595; ROM4[3325]<=26'd23470920;
ROM1[3326]<=26'd1997685; ROM2[3326]<=26'd11312239; ROM3[3326]<=26'd9740939; ROM4[3326]<=26'd23463861;
ROM1[3327]<=26'd1988849; ROM2[3327]<=26'd11311146; ROM3[3327]<=26'd9744944; ROM4[3327]<=26'd23464527;
ROM1[3328]<=26'd1985577; ROM2[3328]<=26'd11312564; ROM3[3328]<=26'd9751045; ROM4[3328]<=26'd23468039;
ROM1[3329]<=26'd1974489; ROM2[3329]<=26'd11308207; ROM3[3329]<=26'd9749635; ROM4[3329]<=26'd23463560;
ROM1[3330]<=26'd1974305; ROM2[3330]<=26'd11309402; ROM3[3330]<=26'd9751169; ROM4[3330]<=26'd23464396;
ROM1[3331]<=26'd1989749; ROM2[3331]<=26'd11319108; ROM3[3331]<=26'd9755313; ROM4[3331]<=26'd23471754;
ROM1[3332]<=26'd2004748; ROM2[3332]<=26'd11322689; ROM3[3332]<=26'd9751459; ROM4[3332]<=26'd23472620;
ROM1[3333]<=26'd2001395; ROM2[3333]<=26'd11312802; ROM3[3333]<=26'd9738716; ROM4[3333]<=26'd23463058;
ROM1[3334]<=26'd1991734; ROM2[3334]<=26'd11307281; ROM3[3334]<=26'd9735809; ROM4[3334]<=26'd23459786;
ROM1[3335]<=26'd1986495; ROM2[3335]<=26'd11308485; ROM3[3335]<=26'd9742779; ROM4[3335]<=26'd23463208;
ROM1[3336]<=26'd1982314; ROM2[3336]<=26'd11310024; ROM3[3336]<=26'd9748197; ROM4[3336]<=26'd23464805;
ROM1[3337]<=26'd1977495; ROM2[3337]<=26'd11311019; ROM3[3337]<=26'd9751471; ROM4[3337]<=26'd23463711;
ROM1[3338]<=26'd1976217; ROM2[3338]<=26'd11312381; ROM3[3338]<=26'd9753855; ROM4[3338]<=26'd23464910;
ROM1[3339]<=26'd1980785; ROM2[3339]<=26'd11313319; ROM3[3339]<=26'd9750956; ROM4[3339]<=26'd23464285;
ROM1[3340]<=26'd1992916; ROM2[3340]<=26'd11314927; ROM3[3340]<=26'd9747882; ROM4[3340]<=26'd23466051;
ROM1[3341]<=26'd2007326; ROM2[3341]<=26'd11320703; ROM3[3341]<=26'd9748541; ROM4[3341]<=26'd23471565;
ROM1[3342]<=26'd2007748; ROM2[3342]<=26'd11323244; ROM3[3342]<=26'd9749744; ROM4[3342]<=26'd23473925;
ROM1[3343]<=26'd2000724; ROM2[3343]<=26'd11321428; ROM3[3343]<=26'd9751180; ROM4[3343]<=26'd23473662;
ROM1[3344]<=26'd1999034; ROM2[3344]<=26'd11322740; ROM3[3344]<=26'd9757611; ROM4[3344]<=26'd23476936;
ROM1[3345]<=26'd1996376; ROM2[3345]<=26'd11323041; ROM3[3345]<=26'd9764637; ROM4[3345]<=26'd23482576;
ROM1[3346]<=26'd1990151; ROM2[3346]<=26'd11322705; ROM3[3346]<=26'd9768599; ROM4[3346]<=26'd23484094;
ROM1[3347]<=26'd1993800; ROM2[3347]<=26'd11325244; ROM3[3347]<=26'd9770555; ROM4[3347]<=26'd23485388;
ROM1[3348]<=26'd2001511; ROM2[3348]<=26'd11323829; ROM3[3348]<=26'd9765871; ROM4[3348]<=26'd23485163;
ROM1[3349]<=26'd2012440; ROM2[3349]<=26'd11323928; ROM3[3349]<=26'd9758565; ROM4[3349]<=26'd23483755;
ROM1[3350]<=26'd2011791; ROM2[3350]<=26'd11322021; ROM3[3350]<=26'd9754337; ROM4[3350]<=26'd23480672;
ROM1[3351]<=26'd1999078; ROM2[3351]<=26'd11317493; ROM3[3351]<=26'd9752888; ROM4[3351]<=26'd23478288;
ROM1[3352]<=26'd1989289; ROM2[3352]<=26'd11316190; ROM3[3352]<=26'd9757571; ROM4[3352]<=26'd23478483;
ROM1[3353]<=26'd1986625; ROM2[3353]<=26'd11316958; ROM3[3353]<=26'd9763307; ROM4[3353]<=26'd23480886;
ROM1[3354]<=26'd1982707; ROM2[3354]<=26'd11316655; ROM3[3354]<=26'd9767378; ROM4[3354]<=26'd23482523;
ROM1[3355]<=26'd1983950; ROM2[3355]<=26'd11317732; ROM3[3355]<=26'd9769578; ROM4[3355]<=26'd23483761;
ROM1[3356]<=26'd1992821; ROM2[3356]<=26'd11321402; ROM3[3356]<=26'd9768312; ROM4[3356]<=26'd23485732;
ROM1[3357]<=26'd2005097; ROM2[3357]<=26'd11323887; ROM3[3357]<=26'd9765378; ROM4[3357]<=26'd23487424;
ROM1[3358]<=26'd2007823; ROM2[3358]<=26'd11321145; ROM3[3358]<=26'd9759575; ROM4[3358]<=26'd23485836;
ROM1[3359]<=26'd2000509; ROM2[3359]<=26'd11317740; ROM3[3359]<=26'd9759887; ROM4[3359]<=26'd23483449;
ROM1[3360]<=26'd1994734; ROM2[3360]<=26'd11319330; ROM3[3360]<=26'd9764109; ROM4[3360]<=26'd23483956;
ROM1[3361]<=26'd1985794; ROM2[3361]<=26'd11316156; ROM3[3361]<=26'd9763352; ROM4[3361]<=26'd23481562;
ROM1[3362]<=26'd1973923; ROM2[3362]<=26'd11309523; ROM3[3362]<=26'd9762934; ROM4[3362]<=26'd23477006;
ROM1[3363]<=26'd1972464; ROM2[3363]<=26'd11309743; ROM3[3363]<=26'd9765483; ROM4[3363]<=26'd23477661;
ROM1[3364]<=26'd1973008; ROM2[3364]<=26'd11305848; ROM3[3364]<=26'd9760136; ROM4[3364]<=26'd23475707;
ROM1[3365]<=26'd1983558; ROM2[3365]<=26'd11305947; ROM3[3365]<=26'd9752882; ROM4[3365]<=26'd23474350;
ROM1[3366]<=26'd2000481; ROM2[3366]<=26'd11313392; ROM3[3366]<=26'd9751938; ROM4[3366]<=26'd23478027;
ROM1[3367]<=26'd1997766; ROM2[3367]<=26'd11310934; ROM3[3367]<=26'd9750974; ROM4[3367]<=26'd23477149;
ROM1[3368]<=26'd1986217; ROM2[3368]<=26'd11306271; ROM3[3368]<=26'd9750833; ROM4[3368]<=26'd23473901;
ROM1[3369]<=26'd1981299; ROM2[3369]<=26'd11307663; ROM3[3369]<=26'd9756860; ROM4[3369]<=26'd23475363;
ROM1[3370]<=26'd1981964; ROM2[3370]<=26'd11313338; ROM3[3370]<=26'd9764813; ROM4[3370]<=26'd23482440;
ROM1[3371]<=26'd1975249; ROM2[3371]<=26'd11311360; ROM3[3371]<=26'd9762966; ROM4[3371]<=26'd23479862;
ROM1[3372]<=26'd1975122; ROM2[3372]<=26'd11309760; ROM3[3372]<=26'd9759517; ROM4[3372]<=26'd23476283;
ROM1[3373]<=26'd1986703; ROM2[3373]<=26'd11314148; ROM3[3373]<=26'd9756883; ROM4[3373]<=26'd23477706;
ROM1[3374]<=26'd2003470; ROM2[3374]<=26'd11317450; ROM3[3374]<=26'd9753685; ROM4[3374]<=26'd23479112;
ROM1[3375]<=26'd2000851; ROM2[3375]<=26'd11314840; ROM3[3375]<=26'd9751813; ROM4[3375]<=26'd23477891;
ROM1[3376]<=26'd1994233; ROM2[3376]<=26'd11314023; ROM3[3376]<=26'd9753181; ROM4[3376]<=26'd23477485;
ROM1[3377]<=26'd1989011; ROM2[3377]<=26'd11312297; ROM3[3377]<=26'd9755015; ROM4[3377]<=26'd23475779;
ROM1[3378]<=26'd1978398; ROM2[3378]<=26'd11307474; ROM3[3378]<=26'd9754186; ROM4[3378]<=26'd23472286;
ROM1[3379]<=26'd1973935; ROM2[3379]<=26'd11307492; ROM3[3379]<=26'd9755924; ROM4[3379]<=26'd23471320;
ROM1[3380]<=26'd1973839; ROM2[3380]<=26'd11308926; ROM3[3380]<=26'd9757790; ROM4[3380]<=26'd23473290;
ROM1[3381]<=26'd1981921; ROM2[3381]<=26'd11313177; ROM3[3381]<=26'd9758901; ROM4[3381]<=26'd23479122;
ROM1[3382]<=26'd1995836; ROM2[3382]<=26'd11314485; ROM3[3382]<=26'd9752656; ROM4[3382]<=26'd23478192;
ROM1[3383]<=26'd2003563; ROM2[3383]<=26'd11315877; ROM3[3383]<=26'd9749972; ROM4[3383]<=26'd23477824;
ROM1[3384]<=26'd2000844; ROM2[3384]<=26'd11317210; ROM3[3384]<=26'd9752388; ROM4[3384]<=26'd23480231;
ROM1[3385]<=26'd1992550; ROM2[3385]<=26'd11315329; ROM3[3385]<=26'd9753226; ROM4[3385]<=26'd23479434;
ROM1[3386]<=26'd1985560; ROM2[3386]<=26'd11315384; ROM3[3386]<=26'd9756587; ROM4[3386]<=26'd23479267;
ROM1[3387]<=26'd1979879; ROM2[3387]<=26'd11316550; ROM3[3387]<=26'd9760938; ROM4[3387]<=26'd23482012;
ROM1[3388]<=26'd1973956; ROM2[3388]<=26'd11313947; ROM3[3388]<=26'd9760493; ROM4[3388]<=26'd23479931;
ROM1[3389]<=26'd1975125; ROM2[3389]<=26'd11310685; ROM3[3389]<=26'd9756303; ROM4[3389]<=26'd23475346;
ROM1[3390]<=26'd1986268; ROM2[3390]<=26'd11312647; ROM3[3390]<=26'd9751102; ROM4[3390]<=26'd23474859;
ROM1[3391]<=26'd1998960; ROM2[3391]<=26'd11317060; ROM3[3391]<=26'd9745832; ROM4[3391]<=26'd23476136;
ROM1[3392]<=26'd1999877; ROM2[3392]<=26'd11319279; ROM3[3392]<=26'd9747310; ROM4[3392]<=26'd23477637;
ROM1[3393]<=26'd1995059; ROM2[3393]<=26'd11320232; ROM3[3393]<=26'd9753182; ROM4[3393]<=26'd23478702;
ROM1[3394]<=26'd1988436; ROM2[3394]<=26'd11320237; ROM3[3394]<=26'd9757036; ROM4[3394]<=26'd23479575;
ROM1[3395]<=26'd1984772; ROM2[3395]<=26'd11322619; ROM3[3395]<=26'd9763274; ROM4[3395]<=26'd23482987;
ROM1[3396]<=26'd1986104; ROM2[3396]<=26'd11328312; ROM3[3396]<=26'd9770305; ROM4[3396]<=26'd23486521;
ROM1[3397]<=26'd1992422; ROM2[3397]<=26'd11332967; ROM3[3397]<=26'd9772940; ROM4[3397]<=26'd23490058;
ROM1[3398]<=26'd2005618; ROM2[3398]<=26'd11335813; ROM3[3398]<=26'd9774442; ROM4[3398]<=26'd23493768;
ROM1[3399]<=26'd2010427; ROM2[3399]<=26'd11327128; ROM3[3399]<=26'd9762546; ROM4[3399]<=26'd23486697;
ROM1[3400]<=26'd2006276; ROM2[3400]<=26'd11319095; ROM3[3400]<=26'd9755129; ROM4[3400]<=26'd23481102;
ROM1[3401]<=26'd2001186; ROM2[3401]<=26'd11320387; ROM3[3401]<=26'd9759750; ROM4[3401]<=26'd23484309;
ROM1[3402]<=26'd1992730; ROM2[3402]<=26'd11319143; ROM3[3402]<=26'd9762738; ROM4[3402]<=26'd23484403;
ROM1[3403]<=26'd1989386; ROM2[3403]<=26'd11317489; ROM3[3403]<=26'd9766581; ROM4[3403]<=26'd23484451;
ROM1[3404]<=26'd1985725; ROM2[3404]<=26'd11318809; ROM3[3404]<=26'd9771753; ROM4[3404]<=26'd23488324;
ROM1[3405]<=26'd1982304; ROM2[3405]<=26'd11314828; ROM3[3405]<=26'd9768246; ROM4[3405]<=26'd23485040;
ROM1[3406]<=26'd1986553; ROM2[3406]<=26'd11312560; ROM3[3406]<=26'd9762459; ROM4[3406]<=26'd23480295;
ROM1[3407]<=26'd2001660; ROM2[3407]<=26'd11317038; ROM3[3407]<=26'd9759131; ROM4[3407]<=26'd23482487;
ROM1[3408]<=26'd2006110; ROM2[3408]<=26'd11316283; ROM3[3408]<=26'd9755142; ROM4[3408]<=26'd23481443;
ROM1[3409]<=26'd1998164; ROM2[3409]<=26'd11313668; ROM3[3409]<=26'd9754770; ROM4[3409]<=26'd23478987;
ROM1[3410]<=26'd1993029; ROM2[3410]<=26'd11312557; ROM3[3410]<=26'd9758740; ROM4[3410]<=26'd23481156;
ROM1[3411]<=26'd1989178; ROM2[3411]<=26'd11314043; ROM3[3411]<=26'd9764049; ROM4[3411]<=26'd23483783;
ROM1[3412]<=26'd1982040; ROM2[3412]<=26'd11314585; ROM3[3412]<=26'd9765767; ROM4[3412]<=26'd23483050;
ROM1[3413]<=26'd1978337; ROM2[3413]<=26'd11314572; ROM3[3413]<=26'd9766436; ROM4[3413]<=26'd23481183;
ROM1[3414]<=26'd1985402; ROM2[3414]<=26'd11318889; ROM3[3414]<=26'd9767472; ROM4[3414]<=26'd23484369;
ROM1[3415]<=26'd2007118; ROM2[3415]<=26'd11331575; ROM3[3415]<=26'd9774072; ROM4[3415]<=26'd23496910;
ROM1[3416]<=26'd2021688; ROM2[3416]<=26'd11334672; ROM3[3416]<=26'd9774418; ROM4[3416]<=26'd23500335;
ROM1[3417]<=26'd2010272; ROM2[3417]<=26'd11322120; ROM3[3417]<=26'd9765614; ROM4[3417]<=26'd23492591;
ROM1[3418]<=26'd2001786; ROM2[3418]<=26'd11319942; ROM3[3418]<=26'd9769211; ROM4[3418]<=26'd23493113;
ROM1[3419]<=26'd1998124; ROM2[3419]<=26'd11322094; ROM3[3419]<=26'd9777055; ROM4[3419]<=26'd23495455;
ROM1[3420]<=26'd1988921; ROM2[3420]<=26'd11317859; ROM3[3420]<=26'd9775741; ROM4[3420]<=26'd23492952;
ROM1[3421]<=26'd1982862; ROM2[3421]<=26'd11314939; ROM3[3421]<=26'd9776168; ROM4[3421]<=26'd23489937;
ROM1[3422]<=26'd1982524; ROM2[3422]<=26'd11312996; ROM3[3422]<=26'd9773537; ROM4[3422]<=26'd23486760;
ROM1[3423]<=26'd1991276; ROM2[3423]<=26'd11311786; ROM3[3423]<=26'd9767843; ROM4[3423]<=26'd23485187;
ROM1[3424]<=26'd2005186; ROM2[3424]<=26'd11313770; ROM3[3424]<=26'd9764068; ROM4[3424]<=26'd23486080;
ROM1[3425]<=26'd2011220; ROM2[3425]<=26'd11316899; ROM3[3425]<=26'd9766112; ROM4[3425]<=26'd23490194;
ROM1[3426]<=26'd2007911; ROM2[3426]<=26'd11318125; ROM3[3426]<=26'd9770805; ROM4[3426]<=26'd23493073;
ROM1[3427]<=26'd1998945; ROM2[3427]<=26'd11317023; ROM3[3427]<=26'd9772571; ROM4[3427]<=26'd23491632;
ROM1[3428]<=26'd1995695; ROM2[3428]<=26'd11318610; ROM3[3428]<=26'd9777549; ROM4[3428]<=26'd23495393;
ROM1[3429]<=26'd1992473; ROM2[3429]<=26'd11319244; ROM3[3429]<=26'd9782423; ROM4[3429]<=26'd23497363;
ROM1[3430]<=26'd1992478; ROM2[3430]<=26'd11319986; ROM3[3430]<=26'd9781027; ROM4[3430]<=26'd23495482;
ROM1[3431]<=26'd1995210; ROM2[3431]<=26'd11317545; ROM3[3431]<=26'd9774149; ROM4[3431]<=26'd23491881;
ROM1[3432]<=26'd2004660; ROM2[3432]<=26'd11316896; ROM3[3432]<=26'd9767023; ROM4[3432]<=26'd23488333;
ROM1[3433]<=26'd2011242; ROM2[3433]<=26'd11321337; ROM3[3433]<=26'd9766075; ROM4[3433]<=26'd23491117;
ROM1[3434]<=26'd2006171; ROM2[3434]<=26'd11320152; ROM3[3434]<=26'd9768323; ROM4[3434]<=26'd23492113;
ROM1[3435]<=26'd1996653; ROM2[3435]<=26'd11317142; ROM3[3435]<=26'd9768860; ROM4[3435]<=26'd23489286;
ROM1[3436]<=26'd1991639; ROM2[3436]<=26'd11318355; ROM3[3436]<=26'd9772232; ROM4[3436]<=26'd23490001;
ROM1[3437]<=26'd1991044; ROM2[3437]<=26'd11322889; ROM3[3437]<=26'd9781284; ROM4[3437]<=26'd23495560;
ROM1[3438]<=26'd1986513; ROM2[3438]<=26'd11321912; ROM3[3438]<=26'd9781678; ROM4[3438]<=26'd23496011;
ROM1[3439]<=26'd1991754; ROM2[3439]<=26'd11321913; ROM3[3439]<=26'd9780329; ROM4[3439]<=26'd23495976;
ROM1[3440]<=26'd2009739; ROM2[3440]<=26'd11326004; ROM3[3440]<=26'd9780160; ROM4[3440]<=26'd23500431;
ROM1[3441]<=26'd2013120; ROM2[3441]<=26'd11319974; ROM3[3441]<=26'd9767317; ROM4[3441]<=26'd23492724;
ROM1[3442]<=26'd2008253; ROM2[3442]<=26'd11317630; ROM3[3442]<=26'd9764198; ROM4[3442]<=26'd23488931;
ROM1[3443]<=26'd2004795; ROM2[3443]<=26'd11318882; ROM3[3443]<=26'd9769376; ROM4[3443]<=26'd23491632;
ROM1[3444]<=26'd1992919; ROM2[3444]<=26'd11312123; ROM3[3444]<=26'd9767648; ROM4[3444]<=26'd23487048;
ROM1[3445]<=26'd1984587; ROM2[3445]<=26'd11311417; ROM3[3445]<=26'd9769026; ROM4[3445]<=26'd23485959;
ROM1[3446]<=26'd1981201; ROM2[3446]<=26'd11313390; ROM3[3446]<=26'd9772546; ROM4[3446]<=26'd23488686;
ROM1[3447]<=26'd1980329; ROM2[3447]<=26'd11311112; ROM3[3447]<=26'd9770638; ROM4[3447]<=26'd23487525;
ROM1[3448]<=26'd1989821; ROM2[3448]<=26'd11310951; ROM3[3448]<=26'd9765198; ROM4[3448]<=26'd23485442;
ROM1[3449]<=26'd2006966; ROM2[3449]<=26'd11316684; ROM3[3449]<=26'd9763892; ROM4[3449]<=26'd23488129;
ROM1[3450]<=26'd2012093; ROM2[3450]<=26'd11319625; ROM3[3450]<=26'd9769284; ROM4[3450]<=26'd23491120;
ROM1[3451]<=26'd2002325; ROM2[3451]<=26'd11316130; ROM3[3451]<=26'd9768806; ROM4[3451]<=26'd23488762;
ROM1[3452]<=26'd1994297; ROM2[3452]<=26'd11317744; ROM3[3452]<=26'd9772065; ROM4[3452]<=26'd23489611;
ROM1[3453]<=26'd1990517; ROM2[3453]<=26'd11318429; ROM3[3453]<=26'd9776148; ROM4[3453]<=26'd23491710;
ROM1[3454]<=26'd1985242; ROM2[3454]<=26'd11319685; ROM3[3454]<=26'd9776931; ROM4[3454]<=26'd23491731;
ROM1[3455]<=26'd1984243; ROM2[3455]<=26'd11319987; ROM3[3455]<=26'd9776660; ROM4[3455]<=26'd23489008;
ROM1[3456]<=26'd1986581; ROM2[3456]<=26'd11315983; ROM3[3456]<=26'd9770134; ROM4[3456]<=26'd23483547;
ROM1[3457]<=26'd2000046; ROM2[3457]<=26'd11318089; ROM3[3457]<=26'd9765498; ROM4[3457]<=26'd23484295;
ROM1[3458]<=26'd2004474; ROM2[3458]<=26'd11316403; ROM3[3458]<=26'd9761894; ROM4[3458]<=26'd23482615;
ROM1[3459]<=26'd1999378; ROM2[3459]<=26'd11316294; ROM3[3459]<=26'd9762075; ROM4[3459]<=26'd23482294;
ROM1[3460]<=26'd1991024; ROM2[3460]<=26'd11316213; ROM3[3460]<=26'd9765550; ROM4[3460]<=26'd23482462;
ROM1[3461]<=26'd1984905; ROM2[3461]<=26'd11313062; ROM3[3461]<=26'd9767066; ROM4[3461]<=26'd23481520;
ROM1[3462]<=26'd1981070; ROM2[3462]<=26'd11311955; ROM3[3462]<=26'd9768961; ROM4[3462]<=26'd23482987;
ROM1[3463]<=26'd1982751; ROM2[3463]<=26'd11314859; ROM3[3463]<=26'd9774157; ROM4[3463]<=26'd23487123;
ROM1[3464]<=26'd1994081; ROM2[3464]<=26'd11321413; ROM3[3464]<=26'd9777488; ROM4[3464]<=26'd23491979;
ROM1[3465]<=26'd2004983; ROM2[3465]<=26'd11321668; ROM3[3465]<=26'd9773270; ROM4[3465]<=26'd23490426;
ROM1[3466]<=26'd2011055; ROM2[3466]<=26'd11318364; ROM3[3466]<=26'd9767745; ROM4[3466]<=26'd23487549;
ROM1[3467]<=26'd2009188; ROM2[3467]<=26'd11320071; ROM3[3467]<=26'd9769072; ROM4[3467]<=26'd23490095;
ROM1[3468]<=26'd2002364; ROM2[3468]<=26'd11319924; ROM3[3468]<=26'd9771701; ROM4[3468]<=26'd23491232;
ROM1[3469]<=26'd1991048; ROM2[3469]<=26'd11314893; ROM3[3469]<=26'd9767974; ROM4[3469]<=26'd23485549;
ROM1[3470]<=26'd1986133; ROM2[3470]<=26'd11314198; ROM3[3470]<=26'd9765156; ROM4[3470]<=26'd23483109;
ROM1[3471]<=26'd1982161; ROM2[3471]<=26'd11312887; ROM3[3471]<=26'd9767023; ROM4[3471]<=26'd23482318;
ROM1[3472]<=26'd1983883; ROM2[3472]<=26'd11312731; ROM3[3472]<=26'd9765899; ROM4[3472]<=26'd23481574;
ROM1[3473]<=26'd1993893; ROM2[3473]<=26'd11315805; ROM3[3473]<=26'd9762908; ROM4[3473]<=26'd23481829;
ROM1[3474]<=26'd2002516; ROM2[3474]<=26'd11315949; ROM3[3474]<=26'd9756737; ROM4[3474]<=26'd23478987;
ROM1[3475]<=26'd2005993; ROM2[3475]<=26'd11319531; ROM3[3475]<=26'd9756808; ROM4[3475]<=26'd23481270;
ROM1[3476]<=26'd1998979; ROM2[3476]<=26'd11317761; ROM3[3476]<=26'd9760127; ROM4[3476]<=26'd23480454;
ROM1[3477]<=26'd1986064; ROM2[3477]<=26'd11311386; ROM3[3477]<=26'd9760236; ROM4[3477]<=26'd23476997;
ROM1[3478]<=26'd1981325; ROM2[3478]<=26'd11310960; ROM3[3478]<=26'd9762687; ROM4[3478]<=26'd23478683;
ROM1[3479]<=26'd1975790; ROM2[3479]<=26'd11308453; ROM3[3479]<=26'd9764616; ROM4[3479]<=26'd23477777;
ROM1[3480]<=26'd1972358; ROM2[3480]<=26'd11305406; ROM3[3480]<=26'd9762583; ROM4[3480]<=26'd23475051;
ROM1[3481]<=26'd1982053; ROM2[3481]<=26'd11309611; ROM3[3481]<=26'd9763194; ROM4[3481]<=26'd23477498;
ROM1[3482]<=26'd1996015; ROM2[3482]<=26'd11312930; ROM3[3482]<=26'd9759898; ROM4[3482]<=26'd23479648;
ROM1[3483]<=26'd2005314; ROM2[3483]<=26'd11318572; ROM3[3483]<=26'd9761416; ROM4[3483]<=26'd23485759;
ROM1[3484]<=26'd2003155; ROM2[3484]<=26'd11320395; ROM3[3484]<=26'd9766540; ROM4[3484]<=26'd23489741;
ROM1[3485]<=26'd2000488; ROM2[3485]<=26'd11322812; ROM3[3485]<=26'd9773083; ROM4[3485]<=26'd23493682;
ROM1[3486]<=26'd1996595; ROM2[3486]<=26'd11324357; ROM3[3486]<=26'd9779542; ROM4[3486]<=26'd23496145;
ROM1[3487]<=26'd1979569; ROM2[3487]<=26'd11312117; ROM3[3487]<=26'd9770263; ROM4[3487]<=26'd23484038;
ROM1[3488]<=26'd1977692; ROM2[3488]<=26'd11311166; ROM3[3488]<=26'd9768561; ROM4[3488]<=26'd23482611;
ROM1[3489]<=26'd1984846; ROM2[3489]<=26'd11313015; ROM3[3489]<=26'd9769381; ROM4[3489]<=26'd23484708;
ROM1[3490]<=26'd1991675; ROM2[3490]<=26'd11310186; ROM3[3490]<=26'd9761139; ROM4[3490]<=26'd23480681;
ROM1[3491]<=26'd2001509; ROM2[3491]<=26'd11311432; ROM3[3491]<=26'd9756042; ROM4[3491]<=26'd23479571;
ROM1[3492]<=26'd1998891; ROM2[3492]<=26'd11310560; ROM3[3492]<=26'd9755229; ROM4[3492]<=26'd23479520;
ROM1[3493]<=26'd1994694; ROM2[3493]<=26'd11313612; ROM3[3493]<=26'd9760532; ROM4[3493]<=26'd23481576;
ROM1[3494]<=26'd1993586; ROM2[3494]<=26'd11316738; ROM3[3494]<=26'd9765816; ROM4[3494]<=26'd23484386;
ROM1[3495]<=26'd1990762; ROM2[3495]<=26'd11317962; ROM3[3495]<=26'd9770343; ROM4[3495]<=26'd23487923;
ROM1[3496]<=26'd1986584; ROM2[3496]<=26'd11319955; ROM3[3496]<=26'd9772768; ROM4[3496]<=26'd23489611;
ROM1[3497]<=26'd1984450; ROM2[3497]<=26'd11317475; ROM3[3497]<=26'd9768582; ROM4[3497]<=26'd23486712;
ROM1[3498]<=26'd1991612; ROM2[3498]<=26'd11316611; ROM3[3498]<=26'd9763953; ROM4[3498]<=26'd23484458;
ROM1[3499]<=26'd2005173; ROM2[3499]<=26'd11320685; ROM3[3499]<=26'd9761116; ROM4[3499]<=26'd23486246;
ROM1[3500]<=26'd2006200; ROM2[3500]<=26'd11321215; ROM3[3500]<=26'd9761176; ROM4[3500]<=26'd23485312;
ROM1[3501]<=26'd1997510; ROM2[3501]<=26'd11316638; ROM3[3501]<=26'd9760643; ROM4[3501]<=26'd23482469;
ROM1[3502]<=26'd1983914; ROM2[3502]<=26'd11308891; ROM3[3502]<=26'd9758127; ROM4[3502]<=26'd23476992;
ROM1[3503]<=26'd1977358; ROM2[3503]<=26'd11306781; ROM3[3503]<=26'd9760428; ROM4[3503]<=26'd23475578;
ROM1[3504]<=26'd1971438; ROM2[3504]<=26'd11307423; ROM3[3504]<=26'd9761474; ROM4[3504]<=26'd23475256;
ROM1[3505]<=26'd1970237; ROM2[3505]<=26'd11309555; ROM3[3505]<=26'd9761178; ROM4[3505]<=26'd23474314;
ROM1[3506]<=26'd1982725; ROM2[3506]<=26'd11314024; ROM3[3506]<=26'd9762756; ROM4[3506]<=26'd23478799;
ROM1[3507]<=26'd1995825; ROM2[3507]<=26'd11314451; ROM3[3507]<=26'd9758921; ROM4[3507]<=26'd23478672;
ROM1[3508]<=26'd2000978; ROM2[3508]<=26'd11313713; ROM3[3508]<=26'd9757585; ROM4[3508]<=26'd23478218;
ROM1[3509]<=26'd1995867; ROM2[3509]<=26'd11314193; ROM3[3509]<=26'd9759966; ROM4[3509]<=26'd23480680;
ROM1[3510]<=26'd1992038; ROM2[3510]<=26'd11319112; ROM3[3510]<=26'd9768166; ROM4[3510]<=26'd23484886;
ROM1[3511]<=26'd1986895; ROM2[3511]<=26'd11317906; ROM3[3511]<=26'd9768781; ROM4[3511]<=26'd23483043;
ROM1[3512]<=26'd1971344; ROM2[3512]<=26'd11306573; ROM3[3512]<=26'd9758573; ROM4[3512]<=26'd23472202;
ROM1[3513]<=26'd1966847; ROM2[3513]<=26'd11303740; ROM3[3513]<=26'd9756397; ROM4[3513]<=26'd23468933;
ROM1[3514]<=26'd1971523; ROM2[3514]<=26'd11304140; ROM3[3514]<=26'd9752637; ROM4[3514]<=26'd23467304;
ROM1[3515]<=26'd1979725; ROM2[3515]<=26'd11304002; ROM3[3515]<=26'd9745210; ROM4[3515]<=26'd23464055;
ROM1[3516]<=26'd1992898; ROM2[3516]<=26'd11308537; ROM3[3516]<=26'd9746129; ROM4[3516]<=26'd23468519;
ROM1[3517]<=26'd1994112; ROM2[3517]<=26'd11310614; ROM3[3517]<=26'd9749256; ROM4[3517]<=26'd23472783;
ROM1[3518]<=26'd1984259; ROM2[3518]<=26'd11306694; ROM3[3518]<=26'd9748971; ROM4[3518]<=26'd23470678;
ROM1[3519]<=26'd1978033; ROM2[3519]<=26'd11304802; ROM3[3519]<=26'd9753207; ROM4[3519]<=26'd23470179;
ROM1[3520]<=26'd1977088; ROM2[3520]<=26'd11309137; ROM3[3520]<=26'd9761061; ROM4[3520]<=26'd23475474;
ROM1[3521]<=26'd1973756; ROM2[3521]<=26'd11308622; ROM3[3521]<=26'd9765456; ROM4[3521]<=26'd23479285;
ROM1[3522]<=26'd1971948; ROM2[3522]<=26'd11304034; ROM3[3522]<=26'd9761740; ROM4[3522]<=26'd23475715;
ROM1[3523]<=26'd1980190; ROM2[3523]<=26'd11304884; ROM3[3523]<=26'd9756266; ROM4[3523]<=26'd23473852;
ROM1[3524]<=26'd1994290; ROM2[3524]<=26'd11307802; ROM3[3524]<=26'd9751895; ROM4[3524]<=26'd23474096;
ROM1[3525]<=26'd1994544; ROM2[3525]<=26'd11305169; ROM3[3525]<=26'd9748842; ROM4[3525]<=26'd23471442;
ROM1[3526]<=26'd1987258; ROM2[3526]<=26'd11303022; ROM3[3526]<=26'd9748949; ROM4[3526]<=26'd23470104;
ROM1[3527]<=26'd1978446; ROM2[3527]<=26'd11299615; ROM3[3527]<=26'd9751088; ROM4[3527]<=26'd23470006;
ROM1[3528]<=26'd1971461; ROM2[3528]<=26'd11295857; ROM3[3528]<=26'd9752340; ROM4[3528]<=26'd23469459;
ROM1[3529]<=26'd1966287; ROM2[3529]<=26'd11295200; ROM3[3529]<=26'd9754916; ROM4[3529]<=26'd23469090;
ROM1[3530]<=26'd1966029; ROM2[3530]<=26'd11296557; ROM3[3530]<=26'd9756023; ROM4[3530]<=26'd23469293;
ROM1[3531]<=26'd1974953; ROM2[3531]<=26'd11299551; ROM3[3531]<=26'd9754357; ROM4[3531]<=26'd23471428;
ROM1[3532]<=26'd1990989; ROM2[3532]<=26'd11304164; ROM3[3532]<=26'd9752172; ROM4[3532]<=26'd23474589;
ROM1[3533]<=26'd2005333; ROM2[3533]<=26'd11312897; ROM3[3533]<=26'd9756398; ROM4[3533]<=26'd23480851;
ROM1[3534]<=26'd2004774; ROM2[3534]<=26'd11315566; ROM3[3534]<=26'd9762289; ROM4[3534]<=26'd23486380;
ROM1[3535]<=26'd1993646; ROM2[3535]<=26'd11309899; ROM3[3535]<=26'd9762027; ROM4[3535]<=26'd23483993;
ROM1[3536]<=26'd1988491; ROM2[3536]<=26'd11310419; ROM3[3536]<=26'd9765582; ROM4[3536]<=26'd23483795;
ROM1[3537]<=26'd1976145; ROM2[3537]<=26'd11306312; ROM3[3537]<=26'd9761602; ROM4[3537]<=26'd23478393;
ROM1[3538]<=26'd1963059; ROM2[3538]<=26'd11296183; ROM3[3538]<=26'd9751429; ROM4[3538]<=26'd23468166;
ROM1[3539]<=26'd1967994; ROM2[3539]<=26'd11299162; ROM3[3539]<=26'd9750857; ROM4[3539]<=26'd23469313;
ROM1[3540]<=26'd1983363; ROM2[3540]<=26'd11304419; ROM3[3540]<=26'd9751139; ROM4[3540]<=26'd23472741;
ROM1[3541]<=26'd1999204; ROM2[3541]<=26'd11311845; ROM3[3541]<=26'd9753872; ROM4[3541]<=26'd23479931;
ROM1[3542]<=26'd1998118; ROM2[3542]<=26'd11313526; ROM3[3542]<=26'd9756259; ROM4[3542]<=26'd23481147;
ROM1[3543]<=26'd1988309; ROM2[3543]<=26'd11309539; ROM3[3543]<=26'd9756779; ROM4[3543]<=26'd23477043;
ROM1[3544]<=26'd1980333; ROM2[3544]<=26'd11305864; ROM3[3544]<=26'd9758518; ROM4[3544]<=26'd23476077;
ROM1[3545]<=26'd1972962; ROM2[3545]<=26'd11303514; ROM3[3545]<=26'd9760092; ROM4[3545]<=26'd23475035;
ROM1[3546]<=26'd1972478; ROM2[3546]<=26'd11307844; ROM3[3546]<=26'd9765682; ROM4[3546]<=26'd23479830;
ROM1[3547]<=26'd1978179; ROM2[3547]<=26'd11310647; ROM3[3547]<=26'd9767579; ROM4[3547]<=26'd23482515;
ROM1[3548]<=26'd1995459; ROM2[3548]<=26'd11318875; ROM3[3548]<=26'd9769393; ROM4[3548]<=26'd23487725;
ROM1[3549]<=26'd2007866; ROM2[3549]<=26'd11320339; ROM3[3549]<=26'd9761973; ROM4[3549]<=26'd23485131;
ROM1[3550]<=26'd2004525; ROM2[3550]<=26'd11316066; ROM3[3550]<=26'd9754618; ROM4[3550]<=26'd23479699;
ROM1[3551]<=26'd1999884; ROM2[3551]<=26'd11319461; ROM3[3551]<=26'd9759036; ROM4[3551]<=26'd23482144;
ROM1[3552]<=26'd1986072; ROM2[3552]<=26'd11313160; ROM3[3552]<=26'd9754468; ROM4[3552]<=26'd23476272;
ROM1[3553]<=26'd1976876; ROM2[3553]<=26'd11307061; ROM3[3553]<=26'd9751450; ROM4[3553]<=26'd23471512;
ROM1[3554]<=26'd1976303; ROM2[3554]<=26'd11312377; ROM3[3554]<=26'd9758588; ROM4[3554]<=26'd23477010;
ROM1[3555]<=26'd1976047; ROM2[3555]<=26'd11311676; ROM3[3555]<=26'd9757008; ROM4[3555]<=26'd23476853;
ROM1[3556]<=26'd1979578; ROM2[3556]<=26'd11309167; ROM3[3556]<=26'd9750242; ROM4[3556]<=26'd23472883;
ROM1[3557]<=26'd1993817; ROM2[3557]<=26'd11312030; ROM3[3557]<=26'd9746212; ROM4[3557]<=26'd23474394;
ROM1[3558]<=26'd2003274; ROM2[3558]<=26'd11315461; ROM3[3558]<=26'd9747832; ROM4[3558]<=26'd23478102;
ROM1[3559]<=26'd1997217; ROM2[3559]<=26'd11313338; ROM3[3559]<=26'd9749866; ROM4[3559]<=26'd23477816;
ROM1[3560]<=26'd1988694; ROM2[3560]<=26'd11309236; ROM3[3560]<=26'd9750976; ROM4[3560]<=26'd23476530;
ROM1[3561]<=26'd1985664; ROM2[3561]<=26'd11311300; ROM3[3561]<=26'd9755289; ROM4[3561]<=26'd23479486;
ROM1[3562]<=26'd1981383; ROM2[3562]<=26'd11312053; ROM3[3562]<=26'd9760367; ROM4[3562]<=26'd23480946;
ROM1[3563]<=26'd1981241; ROM2[3563]<=26'd11314536; ROM3[3563]<=26'd9764903; ROM4[3563]<=26'd23483853;
ROM1[3564]<=26'd1988251; ROM2[3564]<=26'd11321392; ROM3[3564]<=26'd9767883; ROM4[3564]<=26'd23488256;
ROM1[3565]<=26'd1992583; ROM2[3565]<=26'd11314781; ROM3[3565]<=26'd9760344; ROM4[3565]<=26'd23482080;
ROM1[3566]<=26'd1993990; ROM2[3566]<=26'd11305380; ROM3[3566]<=26'd9750693; ROM4[3566]<=26'd23473072;
ROM1[3567]<=26'd1989826; ROM2[3567]<=26'd11303472; ROM3[3567]<=26'd9749884; ROM4[3567]<=26'd23471211;
ROM1[3568]<=26'd1982437; ROM2[3568]<=26'd11301578; ROM3[3568]<=26'd9753651; ROM4[3568]<=26'd23471045;
ROM1[3569]<=26'd1982554; ROM2[3569]<=26'd11305786; ROM3[3569]<=26'd9763979; ROM4[3569]<=26'd23477558;
ROM1[3570]<=26'd1982322; ROM2[3570]<=26'd11309815; ROM3[3570]<=26'd9768767; ROM4[3570]<=26'd23481632;
ROM1[3571]<=26'd1972644; ROM2[3571]<=26'd11304805; ROM3[3571]<=26'd9765052; ROM4[3571]<=26'd23476469;
ROM1[3572]<=26'd1970595; ROM2[3572]<=26'd11299239; ROM3[3572]<=26'd9760920; ROM4[3572]<=26'd23472651;
ROM1[3573]<=26'd1981353; ROM2[3573]<=26'd11301736; ROM3[3573]<=26'd9756905; ROM4[3573]<=26'd23472861;
ROM1[3574]<=26'd1998548; ROM2[3574]<=26'd11308895; ROM3[3574]<=26'd9757126; ROM4[3574]<=26'd23479791;
ROM1[3575]<=26'd2008123; ROM2[3575]<=26'd11316699; ROM3[3575]<=26'd9764196; ROM4[3575]<=26'd23488156;
ROM1[3576]<=26'd1999990; ROM2[3576]<=26'd11313925; ROM3[3576]<=26'd9765027; ROM4[3576]<=26'd23485725;
ROM1[3577]<=26'd1982534; ROM2[3577]<=26'd11304464; ROM3[3577]<=26'd9762586; ROM4[3577]<=26'd23479303;
ROM1[3578]<=26'd1972101; ROM2[3578]<=26'd11299951; ROM3[3578]<=26'd9762270; ROM4[3578]<=26'd23475589;
ROM1[3579]<=26'd1964335; ROM2[3579]<=26'd11296723; ROM3[3579]<=26'd9762048; ROM4[3579]<=26'd23474037;
ROM1[3580]<=26'd1967249; ROM2[3580]<=26'd11300480; ROM3[3580]<=26'd9763870; ROM4[3580]<=26'd23476723;
ROM1[3581]<=26'd1977089; ROM2[3581]<=26'd11303267; ROM3[3581]<=26'd9760852; ROM4[3581]<=26'd23477315;
ROM1[3582]<=26'd1989673; ROM2[3582]<=26'd11302976; ROM3[3582]<=26'd9754840; ROM4[3582]<=26'd23477060;
ROM1[3583]<=26'd1995260; ROM2[3583]<=26'd11305377; ROM3[3583]<=26'd9753154; ROM4[3583]<=26'd23477883;
ROM1[3584]<=26'd1990919; ROM2[3584]<=26'd11307397; ROM3[3584]<=26'd9756100; ROM4[3584]<=26'd23479091;
ROM1[3585]<=26'd1986541; ROM2[3585]<=26'd11310381; ROM3[3585]<=26'd9760693; ROM4[3585]<=26'd23481438;
ROM1[3586]<=26'd1984547; ROM2[3586]<=26'd11313694; ROM3[3586]<=26'd9764995; ROM4[3586]<=26'd23483266;
ROM1[3587]<=26'd1978679; ROM2[3587]<=26'd11310097; ROM3[3587]<=26'd9764602; ROM4[3587]<=26'd23480461;
ROM1[3588]<=26'd1974809; ROM2[3588]<=26'd11306912; ROM3[3588]<=26'd9763439; ROM4[3588]<=26'd23478994;
ROM1[3589]<=26'd1975879; ROM2[3589]<=26'd11305966; ROM3[3589]<=26'd9759949; ROM4[3589]<=26'd23475314;
ROM1[3590]<=26'd1985723; ROM2[3590]<=26'd11305404; ROM3[3590]<=26'd9752397; ROM4[3590]<=26'd23472202;
ROM1[3591]<=26'd1994860; ROM2[3591]<=26'd11305085; ROM3[3591]<=26'd9746136; ROM4[3591]<=26'd23470621;
ROM1[3592]<=26'd1991777; ROM2[3592]<=26'd11303853; ROM3[3592]<=26'd9745134; ROM4[3592]<=26'd23467768;
ROM1[3593]<=26'd1991508; ROM2[3593]<=26'd11308593; ROM3[3593]<=26'd9752847; ROM4[3593]<=26'd23472336;
ROM1[3594]<=26'd1994417; ROM2[3594]<=26'd11316928; ROM3[3594]<=26'd9765274; ROM4[3594]<=26'd23480224;
ROM1[3595]<=26'd1989285; ROM2[3595]<=26'd11315325; ROM3[3595]<=26'd9767449; ROM4[3595]<=26'd23479246;
ROM1[3596]<=26'd1976717; ROM2[3596]<=26'd11306248; ROM3[3596]<=26'd9759076; ROM4[3596]<=26'd23469293;
ROM1[3597]<=26'd1977331; ROM2[3597]<=26'd11304888; ROM3[3597]<=26'd9755145; ROM4[3597]<=26'd23466882;
ROM1[3598]<=26'd1987473; ROM2[3598]<=26'd11306533; ROM3[3598]<=26'd9752269; ROM4[3598]<=26'd23467296;
ROM1[3599]<=26'd1999960; ROM2[3599]<=26'd11311637; ROM3[3599]<=26'd9747867; ROM4[3599]<=26'd23467160;
ROM1[3600]<=26'd2005918; ROM2[3600]<=26'd11317292; ROM3[3600]<=26'd9751516; ROM4[3600]<=26'd23472835;
ROM1[3601]<=26'd1998197; ROM2[3601]<=26'd11316276; ROM3[3601]<=26'd9755387; ROM4[3601]<=26'd23474221;
ROM1[3602]<=26'd1985003; ROM2[3602]<=26'd11310784; ROM3[3602]<=26'd9755458; ROM4[3602]<=26'd23471688;
ROM1[3603]<=26'd1979442; ROM2[3603]<=26'd11309317; ROM3[3603]<=26'd9760912; ROM4[3603]<=26'd23473397;
ROM1[3604]<=26'd1976221; ROM2[3604]<=26'd11311369; ROM3[3604]<=26'd9768360; ROM4[3604]<=26'd23477104;
ROM1[3605]<=26'd1976520; ROM2[3605]<=26'd11311258; ROM3[3605]<=26'd9769782; ROM4[3605]<=26'd23476518;
ROM1[3606]<=26'd1979160; ROM2[3606]<=26'd11306077; ROM3[3606]<=26'd9761424; ROM4[3606]<=26'd23470014;
ROM1[3607]<=26'd1991115; ROM2[3607]<=26'd11304417; ROM3[3607]<=26'd9754789; ROM4[3607]<=26'd23468786;
ROM1[3608]<=26'd1998791; ROM2[3608]<=26'd11306873; ROM3[3608]<=26'd9756054; ROM4[3608]<=26'd23472549;
ROM1[3609]<=26'd1993119; ROM2[3609]<=26'd11306081; ROM3[3609]<=26'd9759023; ROM4[3609]<=26'd23475211;
ROM1[3610]<=26'd1987899; ROM2[3610]<=26'd11305977; ROM3[3610]<=26'd9763570; ROM4[3610]<=26'd23476367;
ROM1[3611]<=26'd1986022; ROM2[3611]<=26'd11307776; ROM3[3611]<=26'd9769743; ROM4[3611]<=26'd23478870;
ROM1[3612]<=26'd1984331; ROM2[3612]<=26'd11309757; ROM3[3612]<=26'd9773562; ROM4[3612]<=26'd23482081;
ROM1[3613]<=26'd1982211; ROM2[3613]<=26'd11309566; ROM3[3613]<=26'd9773009; ROM4[3613]<=26'd23481901;
ROM1[3614]<=26'd1988111; ROM2[3614]<=26'd11312409; ROM3[3614]<=26'd9772945; ROM4[3614]<=26'd23484021;
ROM1[3615]<=26'd2000489; ROM2[3615]<=26'd11314432; ROM3[3615]<=26'd9768668; ROM4[3615]<=26'd23485954;
ROM1[3616]<=26'd2008859; ROM2[3616]<=26'd11313080; ROM3[3616]<=26'd9763986; ROM4[3616]<=26'd23485600;
ROM1[3617]<=26'd2010846; ROM2[3617]<=26'd11317037; ROM3[3617]<=26'd9769374; ROM4[3617]<=26'd23491094;
ROM1[3618]<=26'd2003023; ROM2[3618]<=26'd11314759; ROM3[3618]<=26'd9772542; ROM4[3618]<=26'd23491661;
ROM1[3619]<=26'd1989972; ROM2[3619]<=26'd11307283; ROM3[3619]<=26'd9771050; ROM4[3619]<=26'd23487181;
ROM1[3620]<=26'd1980751; ROM2[3620]<=26'd11302404; ROM3[3620]<=26'd9770120; ROM4[3620]<=26'd23485393;
ROM1[3621]<=26'd1971700; ROM2[3621]<=26'd11295583; ROM3[3621]<=26'd9766408; ROM4[3621]<=26'd23479182;
ROM1[3622]<=26'd1975343; ROM2[3622]<=26'd11297377; ROM3[3622]<=26'd9765929; ROM4[3622]<=26'd23479400;
ROM1[3623]<=26'd1986465; ROM2[3623]<=26'd11300469; ROM3[3623]<=26'd9765221; ROM4[3623]<=26'd23480384;
ROM1[3624]<=26'd1999194; ROM2[3624]<=26'd11301108; ROM3[3624]<=26'd9761341; ROM4[3624]<=26'd23479595;
ROM1[3625]<=26'd1999507; ROM2[3625]<=26'd11297808; ROM3[3625]<=26'd9758168; ROM4[3625]<=26'd23477960;
ROM1[3626]<=26'd1990607; ROM2[3626]<=26'd11294500; ROM3[3626]<=26'd9757772; ROM4[3626]<=26'd23475539;
ROM1[3627]<=26'd1991710; ROM2[3627]<=26'd11303396; ROM3[3627]<=26'd9768058; ROM4[3627]<=26'd23483338;
ROM1[3628]<=26'd1989178; ROM2[3628]<=26'd11306186; ROM3[3628]<=26'd9771466; ROM4[3628]<=26'd23485465;
ROM1[3629]<=26'd1971085; ROM2[3629]<=26'd11293476; ROM3[3629]<=26'd9762830; ROM4[3629]<=26'd23472221;
ROM1[3630]<=26'd1965542; ROM2[3630]<=26'd11290984; ROM3[3630]<=26'd9759093; ROM4[3630]<=26'd23466991;
ROM1[3631]<=26'd1971528; ROM2[3631]<=26'd11291794; ROM3[3631]<=26'd9753110; ROM4[3631]<=26'd23463896;
ROM1[3632]<=26'd1986499; ROM2[3632]<=26'd11295292; ROM3[3632]<=26'd9747890; ROM4[3632]<=26'd23463024;
ROM1[3633]<=26'd2001774; ROM2[3633]<=26'd11306512; ROM3[3633]<=26'd9750139; ROM4[3633]<=26'd23470567;
ROM1[3634]<=26'd2003521; ROM2[3634]<=26'd11311601; ROM3[3634]<=26'd9755841; ROM4[3634]<=26'd23475920;
ROM1[3635]<=26'd1997003; ROM2[3635]<=26'd11311620; ROM3[3635]<=26'd9760565; ROM4[3635]<=26'd23477535;
ROM1[3636]<=26'd1989734; ROM2[3636]<=26'd11311302; ROM3[3636]<=26'd9762092; ROM4[3636]<=26'd23476733;
ROM1[3637]<=26'd1979773; ROM2[3637]<=26'd11308457; ROM3[3637]<=26'd9762558; ROM4[3637]<=26'd23474720;
ROM1[3638]<=26'd1975425; ROM2[3638]<=26'd11306837; ROM3[3638]<=26'd9761438; ROM4[3638]<=26'd23473598;
ROM1[3639]<=26'd1981419; ROM2[3639]<=26'd11308163; ROM3[3639]<=26'd9758487; ROM4[3639]<=26'd23472475;
ROM1[3640]<=26'd1991248; ROM2[3640]<=26'd11308369; ROM3[3640]<=26'd9751106; ROM4[3640]<=26'd23469910;
ROM1[3641]<=26'd2003345; ROM2[3641]<=26'd11312425; ROM3[3641]<=26'd9750102; ROM4[3641]<=26'd23473149;
ROM1[3642]<=26'd1999970; ROM2[3642]<=26'd11311061; ROM3[3642]<=26'd9750914; ROM4[3642]<=26'd23472588;
ROM1[3643]<=26'd1988071; ROM2[3643]<=26'd11304969; ROM3[3643]<=26'd9749359; ROM4[3643]<=26'd23467750;
ROM1[3644]<=26'd1980096; ROM2[3644]<=26'd11303449; ROM3[3644]<=26'd9752359; ROM4[3644]<=26'd23466585;
ROM1[3645]<=26'd1976920; ROM2[3645]<=26'd11304771; ROM3[3645]<=26'd9755290; ROM4[3645]<=26'd23467808;
ROM1[3646]<=26'd1972140; ROM2[3646]<=26'd11305387; ROM3[3646]<=26'd9756069; ROM4[3646]<=26'd23466822;
ROM1[3647]<=26'd1972169; ROM2[3647]<=26'd11302960; ROM3[3647]<=26'd9751847; ROM4[3647]<=26'd23463949;
ROM1[3648]<=26'd1981701; ROM2[3648]<=26'd11300331; ROM3[3648]<=26'd9747291; ROM4[3648]<=26'd23461423;
ROM1[3649]<=26'd1995678; ROM2[3649]<=26'd11302905; ROM3[3649]<=26'd9744241; ROM4[3649]<=26'd23461822;
ROM1[3650]<=26'd2000086; ROM2[3650]<=26'd11305991; ROM3[3650]<=26'd9744836; ROM4[3650]<=26'd23464114;
ROM1[3651]<=26'd1991623; ROM2[3651]<=26'd11303884; ROM3[3651]<=26'd9745428; ROM4[3651]<=26'd23462192;
ROM1[3652]<=26'd1983318; ROM2[3652]<=26'd11302349; ROM3[3652]<=26'd9746381; ROM4[3652]<=26'd23461129;
ROM1[3653]<=26'd1981749; ROM2[3653]<=26'd11305220; ROM3[3653]<=26'd9751785; ROM4[3653]<=26'd23464807;
ROM1[3654]<=26'd1978334; ROM2[3654]<=26'd11306343; ROM3[3654]<=26'd9755153; ROM4[3654]<=26'd23465923;
ROM1[3655]<=26'd1977886; ROM2[3655]<=26'd11305189; ROM3[3655]<=26'd9755147; ROM4[3655]<=26'd23465339;
ROM1[3656]<=26'd1986517; ROM2[3656]<=26'd11307875; ROM3[3656]<=26'd9753622; ROM4[3656]<=26'd23466906;
ROM1[3657]<=26'd1996810; ROM2[3657]<=26'd11307042; ROM3[3657]<=26'd9746043; ROM4[3657]<=26'd23465464;
ROM1[3658]<=26'd1998948; ROM2[3658]<=26'd11302162; ROM3[3658]<=26'd9743249; ROM4[3658]<=26'd23463706;
ROM1[3659]<=26'd1997460; ROM2[3659]<=26'd11305430; ROM3[3659]<=26'd9747330; ROM4[3659]<=26'd23467327;
ROM1[3660]<=26'd1995189; ROM2[3660]<=26'd11310777; ROM3[3660]<=26'd9753562; ROM4[3660]<=26'd23473187;
ROM1[3661]<=26'd1991825; ROM2[3661]<=26'd11309101; ROM3[3661]<=26'd9756109; ROM4[3661]<=26'd23472302;
ROM1[3662]<=26'd1984548; ROM2[3662]<=26'd11307205; ROM3[3662]<=26'd9755146; ROM4[3662]<=26'd23468981;
ROM1[3663]<=26'd1985582; ROM2[3663]<=26'd11311697; ROM3[3663]<=26'd9760177; ROM4[3663]<=26'd23474445;
ROM1[3664]<=26'd1996781; ROM2[3664]<=26'd11318116; ROM3[3664]<=26'd9764731; ROM4[3664]<=26'd23481832;
ROM1[3665]<=26'd2011431; ROM2[3665]<=26'd11322984; ROM3[3665]<=26'd9762424; ROM4[3665]<=26'd23484708;
ROM1[3666]<=26'd2017388; ROM2[3666]<=26'd11320324; ROM3[3666]<=26'd9753637; ROM4[3666]<=26'd23480386;
ROM1[3667]<=26'd2007709; ROM2[3667]<=26'd11313160; ROM3[3667]<=26'd9748429; ROM4[3667]<=26'd23474322;
ROM1[3668]<=26'd1993897; ROM2[3668]<=26'd11305765; ROM3[3668]<=26'd9746721; ROM4[3668]<=26'd23469595;
ROM1[3669]<=26'd1983436; ROM2[3669]<=26'd11302611; ROM3[3669]<=26'd9747112; ROM4[3669]<=26'd23467867;
ROM1[3670]<=26'd1985295; ROM2[3670]<=26'd11309589; ROM3[3670]<=26'd9757344; ROM4[3670]<=26'd23476088;
ROM1[3671]<=26'd1990220; ROM2[3671]<=26'd11316472; ROM3[3671]<=26'd9768029; ROM4[3671]<=26'd23484090;
ROM1[3672]<=26'd1986373; ROM2[3672]<=26'd11310110; ROM3[3672]<=26'd9762260; ROM4[3672]<=26'd23478687;
ROM1[3673]<=26'd1995078; ROM2[3673]<=26'd11309720; ROM3[3673]<=26'd9757929; ROM4[3673]<=26'd23476859;
ROM1[3674]<=26'd2006417; ROM2[3674]<=26'd11309746; ROM3[3674]<=26'd9752110; ROM4[3674]<=26'd23477050;
ROM1[3675]<=26'd1997792; ROM2[3675]<=26'd11301607; ROM3[3675]<=26'd9743347; ROM4[3675]<=26'd23470302;
ROM1[3676]<=26'd1993587; ROM2[3676]<=26'd11303537; ROM3[3676]<=26'd9750512; ROM4[3676]<=26'd23472328;
ROM1[3677]<=26'd1988974; ROM2[3677]<=26'd11304967; ROM3[3677]<=26'd9759218; ROM4[3677]<=26'd23476640;
ROM1[3678]<=26'd1984584; ROM2[3678]<=26'd11304848; ROM3[3678]<=26'd9764169; ROM4[3678]<=26'd23478125;
ROM1[3679]<=26'd1982474; ROM2[3679]<=26'd11306650; ROM3[3679]<=26'd9769804; ROM4[3679]<=26'd23481333;
ROM1[3680]<=26'd1982553; ROM2[3680]<=26'd11307264; ROM3[3680]<=26'd9769927; ROM4[3680]<=26'd23481871;
ROM1[3681]<=26'd1987597; ROM2[3681]<=26'd11306127; ROM3[3681]<=26'd9765157; ROM4[3681]<=26'd23479122;
ROM1[3682]<=26'd2002667; ROM2[3682]<=26'd11310050; ROM3[3682]<=26'd9763795; ROM4[3682]<=26'd23481703;
ROM1[3683]<=26'd2011753; ROM2[3683]<=26'd11314876; ROM3[3683]<=26'd9763915; ROM4[3683]<=26'd23484067;
ROM1[3684]<=26'd2000717; ROM2[3684]<=26'd11309269; ROM3[3684]<=26'd9760159; ROM4[3684]<=26'd23477125;
ROM1[3685]<=26'd1984467; ROM2[3685]<=26'd11300524; ROM3[3685]<=26'd9757145; ROM4[3685]<=26'd23471027;
ROM1[3686]<=26'd1973335; ROM2[3686]<=26'd11294830; ROM3[3686]<=26'd9755335; ROM4[3686]<=26'd23466598;
ROM1[3687]<=26'd1961050; ROM2[3687]<=26'd11288571; ROM3[3687]<=26'd9752139; ROM4[3687]<=26'd23459618;
ROM1[3688]<=26'd1958690; ROM2[3688]<=26'd11288918; ROM3[3688]<=26'd9749950; ROM4[3688]<=26'd23458400;
ROM1[3689]<=26'd1966740; ROM2[3689]<=26'd11292826; ROM3[3689]<=26'd9748063; ROM4[3689]<=26'd23460563;
ROM1[3690]<=26'd1978461; ROM2[3690]<=26'd11293752; ROM3[3690]<=26'd9742773; ROM4[3690]<=26'd23459951;
ROM1[3691]<=26'd1989363; ROM2[3691]<=26'd11297842; ROM3[3691]<=26'd9741104; ROM4[3691]<=26'd23462858;
ROM1[3692]<=26'd1988944; ROM2[3692]<=26'd11298854; ROM3[3692]<=26'd9743945; ROM4[3692]<=26'd23466832;
ROM1[3693]<=26'd1981954; ROM2[3693]<=26'd11298094; ROM3[3693]<=26'd9745630; ROM4[3693]<=26'd23466213;
ROM1[3694]<=26'd1975222; ROM2[3694]<=26'd11298780; ROM3[3694]<=26'd9747316; ROM4[3694]<=26'd23464795;
ROM1[3695]<=26'd1969278; ROM2[3695]<=26'd11295376; ROM3[3695]<=26'd9746587; ROM4[3695]<=26'd23463966;
ROM1[3696]<=26'd1968097; ROM2[3696]<=26'd11295929; ROM3[3696]<=26'd9748678; ROM4[3696]<=26'd23466157;
ROM1[3697]<=26'd1974023; ROM2[3697]<=26'd11299020; ROM3[3697]<=26'd9749439; ROM4[3697]<=26'd23467789;
ROM1[3698]<=26'd1986629; ROM2[3698]<=26'd11302635; ROM3[3698]<=26'd9745611; ROM4[3698]<=26'd23469610;
ROM1[3699]<=26'd1999319; ROM2[3699]<=26'd11305596; ROM3[3699]<=26'd9739857; ROM4[3699]<=26'd23469112;
ROM1[3700]<=26'd2001642; ROM2[3700]<=26'd11308845; ROM3[3700]<=26'd9741685; ROM4[3700]<=26'd23469664;
ROM1[3701]<=26'd2003336; ROM2[3701]<=26'd11315701; ROM3[3701]<=26'd9751979; ROM4[3701]<=26'd23477328;
ROM1[3702]<=26'd1995807; ROM2[3702]<=26'd11313381; ROM3[3702]<=26'd9752696; ROM4[3702]<=26'd23476093;
ROM1[3703]<=26'd1984882; ROM2[3703]<=26'd11307724; ROM3[3703]<=26'd9748277; ROM4[3703]<=26'd23469466;
ROM1[3704]<=26'd1976517; ROM2[3704]<=26'd11307205; ROM3[3704]<=26'd9748316; ROM4[3704]<=26'd23468430;
ROM1[3705]<=26'd1973309; ROM2[3705]<=26'd11305368; ROM3[3705]<=26'd9744886; ROM4[3705]<=26'd23466684;
ROM1[3706]<=26'd1981693; ROM2[3706]<=26'd11304783; ROM3[3706]<=26'd9741690; ROM4[3706]<=26'd23465042;
ROM1[3707]<=26'd2000130; ROM2[3707]<=26'd11310180; ROM3[3707]<=26'd9740680; ROM4[3707]<=26'd23469014;
ROM1[3708]<=26'd2009338; ROM2[3708]<=26'd11312551; ROM3[3708]<=26'd9741865; ROM4[3708]<=26'd23473384;
ROM1[3709]<=26'd2005094; ROM2[3709]<=26'd11312023; ROM3[3709]<=26'd9746303; ROM4[3709]<=26'd23473984;
ROM1[3710]<=26'd1993009; ROM2[3710]<=26'd11307085; ROM3[3710]<=26'd9747218; ROM4[3710]<=26'd23471111;
ROM1[3711]<=26'd1986082; ROM2[3711]<=26'd11305880; ROM3[3711]<=26'd9751476; ROM4[3711]<=26'd23472349;
ROM1[3712]<=26'd1982772; ROM2[3712]<=26'd11307182; ROM3[3712]<=26'd9756598; ROM4[3712]<=26'd23473808;
ROM1[3713]<=26'd1979630; ROM2[3713]<=26'd11304891; ROM3[3713]<=26'd9753702; ROM4[3713]<=26'd23469286;
ROM1[3714]<=26'd1989841; ROM2[3714]<=26'd11312943; ROM3[3714]<=26'd9756264; ROM4[3714]<=26'd23472229;
ROM1[3715]<=26'd2007226; ROM2[3715]<=26'd11320236; ROM3[3715]<=26'd9757259; ROM4[3715]<=26'd23478328;
ROM1[3716]<=26'd2008675; ROM2[3716]<=26'd11312957; ROM3[3716]<=26'd9745017; ROM4[3716]<=26'd23470080;
ROM1[3717]<=26'd2002858; ROM2[3717]<=26'd11309280; ROM3[3717]<=26'd9743507; ROM4[3717]<=26'd23468197;
ROM1[3718]<=26'd2001131; ROM2[3718]<=26'd11313519; ROM3[3718]<=26'd9752564; ROM4[3718]<=26'd23476965;
ROM1[3719]<=26'd1992349; ROM2[3719]<=26'd11310408; ROM3[3719]<=26'd9753771; ROM4[3719]<=26'd23475158;
ROM1[3720]<=26'd1987546; ROM2[3720]<=26'd11310852; ROM3[3720]<=26'd9756638; ROM4[3720]<=26'd23474881;
ROM1[3721]<=26'd1981363; ROM2[3721]<=26'd11310984; ROM3[3721]<=26'd9760008; ROM4[3721]<=26'd23474843;
ROM1[3722]<=26'd1977957; ROM2[3722]<=26'd11306588; ROM3[3722]<=26'd9754144; ROM4[3722]<=26'd23470506;
ROM1[3723]<=26'd1989888; ROM2[3723]<=26'd11308505; ROM3[3723]<=26'd9751885; ROM4[3723]<=26'd23471482;
ROM1[3724]<=26'd2003205; ROM2[3724]<=26'd11311261; ROM3[3724]<=26'd9750617; ROM4[3724]<=26'd23472620;
ROM1[3725]<=26'd2003346; ROM2[3725]<=26'd11310554; ROM3[3725]<=26'd9748781; ROM4[3725]<=26'd23471747;
ROM1[3726]<=26'd2000438; ROM2[3726]<=26'd11312228; ROM3[3726]<=26'd9756147; ROM4[3726]<=26'd23475491;
ROM1[3727]<=26'd1998705; ROM2[3727]<=26'd11316758; ROM3[3727]<=26'd9765499; ROM4[3727]<=26'd23480461;
ROM1[3728]<=26'd1993752; ROM2[3728]<=26'd11315379; ROM3[3728]<=26'd9766571; ROM4[3728]<=26'd23481866;
ROM1[3729]<=26'd1980565; ROM2[3729]<=26'd11306578; ROM3[3729]<=26'd9762487; ROM4[3729]<=26'd23474643;
ROM1[3730]<=26'd1974964; ROM2[3730]<=26'd11301624; ROM3[3730]<=26'd9758045; ROM4[3730]<=26'd23469266;
ROM1[3731]<=26'd1977682; ROM2[3731]<=26'd11297613; ROM3[3731]<=26'd9749837; ROM4[3731]<=26'd23465448;
ROM1[3732]<=26'd1991709; ROM2[3732]<=26'd11301428; ROM3[3732]<=26'd9745420; ROM4[3732]<=26'd23464354;
ROM1[3733]<=26'd2001893; ROM2[3733]<=26'd11306684; ROM3[3733]<=26'd9745940; ROM4[3733]<=26'd23469056;
ROM1[3734]<=26'd1995890; ROM2[3734]<=26'd11304758; ROM3[3734]<=26'd9746413; ROM4[3734]<=26'd23468603;
ROM1[3735]<=26'd1987357; ROM2[3735]<=26'd11301518; ROM3[3735]<=26'd9748949; ROM4[3735]<=26'd23466928;
ROM1[3736]<=26'd1988860; ROM2[3736]<=26'd11305701; ROM3[3736]<=26'd9758831; ROM4[3736]<=26'd23474243;
ROM1[3737]<=26'd1988484; ROM2[3737]<=26'd11309810; ROM3[3737]<=26'd9766423; ROM4[3737]<=26'd23479629;
ROM1[3738]<=26'd1983273; ROM2[3738]<=26'd11305334; ROM3[3738]<=26'd9762296; ROM4[3738]<=26'd23475522;
ROM1[3739]<=26'd1987802; ROM2[3739]<=26'd11305157; ROM3[3739]<=26'd9758406; ROM4[3739]<=26'd23472915;
ROM1[3740]<=26'd1997302; ROM2[3740]<=26'd11303572; ROM3[3740]<=26'd9750701; ROM4[3740]<=26'd23469338;
ROM1[3741]<=26'd2005230; ROM2[3741]<=26'd11303870; ROM3[3741]<=26'd9744728; ROM4[3741]<=26'd23469278;
ROM1[3742]<=26'd2004759; ROM2[3742]<=26'd11304876; ROM3[3742]<=26'd9747814; ROM4[3742]<=26'd23471143;
ROM1[3743]<=26'd1995945; ROM2[3743]<=26'd11302073; ROM3[3743]<=26'd9748509; ROM4[3743]<=26'd23469353;
ROM1[3744]<=26'd1987165; ROM2[3744]<=26'd11300712; ROM3[3744]<=26'd9748884; ROM4[3744]<=26'd23468262;
ROM1[3745]<=26'd1986847; ROM2[3745]<=26'd11305282; ROM3[3745]<=26'd9755731; ROM4[3745]<=26'd23472928;
ROM1[3746]<=26'd1985818; ROM2[3746]<=26'd11311310; ROM3[3746]<=26'd9761694; ROM4[3746]<=26'd23477842;
ROM1[3747]<=26'd1981049; ROM2[3747]<=26'd11306394; ROM3[3747]<=26'd9755822; ROM4[3747]<=26'd23472528;
ROM1[3748]<=26'd1986093; ROM2[3748]<=26'd11300549; ROM3[3748]<=26'd9746983; ROM4[3748]<=26'd23466776;
ROM1[3749]<=26'd1999676; ROM2[3749]<=26'd11303637; ROM3[3749]<=26'd9743710; ROM4[3749]<=26'd23468784;
ROM1[3750]<=26'd2001509; ROM2[3750]<=26'd11306170; ROM3[3750]<=26'd9744145; ROM4[3750]<=26'd23471181;
ROM1[3751]<=26'd1990553; ROM2[3751]<=26'd11301401; ROM3[3751]<=26'd9741476; ROM4[3751]<=26'd23467211;
ROM1[3752]<=26'd1975972; ROM2[3752]<=26'd11296322; ROM3[3752]<=26'd9740163; ROM4[3752]<=26'd23463530;
ROM1[3753]<=26'd1966828; ROM2[3753]<=26'd11293233; ROM3[3753]<=26'd9740422; ROM4[3753]<=26'd23460871;
ROM1[3754]<=26'd1959232; ROM2[3754]<=26'd11289135; ROM3[3754]<=26'd9740094; ROM4[3754]<=26'd23458299;
ROM1[3755]<=26'd1965247; ROM2[3755]<=26'd11295447; ROM3[3755]<=26'd9747301; ROM4[3755]<=26'd23464577;
ROM1[3756]<=26'd1977436; ROM2[3756]<=26'd11301582; ROM3[3756]<=26'd9749296; ROM4[3756]<=26'd23469925;
ROM1[3757]<=26'd1988582; ROM2[3757]<=26'd11301401; ROM3[3757]<=26'd9742307; ROM4[3757]<=26'd23468270;
ROM1[3758]<=26'd1993414; ROM2[3758]<=26'd11301205; ROM3[3758]<=26'd9739420; ROM4[3758]<=26'd23467310;
ROM1[3759]<=26'd1992645; ROM2[3759]<=26'd11304185; ROM3[3759]<=26'd9745206; ROM4[3759]<=26'd23472112;
ROM1[3760]<=26'd1988142; ROM2[3760]<=26'd11303938; ROM3[3760]<=26'd9751118; ROM4[3760]<=26'd23473698;
ROM1[3761]<=26'd1982269; ROM2[3761]<=26'd11301197; ROM3[3761]<=26'd9752258; ROM4[3761]<=26'd23472002;
ROM1[3762]<=26'd1975987; ROM2[3762]<=26'd11300435; ROM3[3762]<=26'd9753861; ROM4[3762]<=26'd23471663;
ROM1[3763]<=26'd1975134; ROM2[3763]<=26'd11300700; ROM3[3763]<=26'd9758472; ROM4[3763]<=26'd23473272;
ROM1[3764]<=26'd1979411; ROM2[3764]<=26'd11301341; ROM3[3764]<=26'd9756317; ROM4[3764]<=26'd23471928;
ROM1[3765]<=26'd1989820; ROM2[3765]<=26'd11301533; ROM3[3765]<=26'd9748396; ROM4[3765]<=26'd23470422;
ROM1[3766]<=26'd1998204; ROM2[3766]<=26'd11299973; ROM3[3766]<=26'd9742095; ROM4[3766]<=26'd23468493;
ROM1[3767]<=26'd1997372; ROM2[3767]<=26'd11300948; ROM3[3767]<=26'd9742143; ROM4[3767]<=26'd23467285;
ROM1[3768]<=26'd1995599; ROM2[3768]<=26'd11303145; ROM3[3768]<=26'd9749853; ROM4[3768]<=26'd23473091;
ROM1[3769]<=26'd1991953; ROM2[3769]<=26'd11304455; ROM3[3769]<=26'd9757580; ROM4[3769]<=26'd23476576;
ROM1[3770]<=26'd1994403; ROM2[3770]<=26'd11311019; ROM3[3770]<=26'd9767892; ROM4[3770]<=26'd23484208;
ROM1[3771]<=26'd1994459; ROM2[3771]<=26'd11314537; ROM3[3771]<=26'd9772093; ROM4[3771]<=26'd23488032;
ROM1[3772]<=26'd1991143; ROM2[3772]<=26'd11309938; ROM3[3772]<=26'd9765307; ROM4[3772]<=26'd23480259;
ROM1[3773]<=26'd1992507; ROM2[3773]<=26'd11303051; ROM3[3773]<=26'd9754137; ROM4[3773]<=26'd23471515;
ROM1[3774]<=26'd1999299; ROM2[3774]<=26'd11300071; ROM3[3774]<=26'd9745232; ROM4[3774]<=26'd23465989;
ROM1[3775]<=26'd1998318; ROM2[3775]<=26'd11298429; ROM3[3775]<=26'd9743093; ROM4[3775]<=26'd23464967;
ROM1[3776]<=26'd1991809; ROM2[3776]<=26'd11299523; ROM3[3776]<=26'd9745562; ROM4[3776]<=26'd23466036;
ROM1[3777]<=26'd1990892; ROM2[3777]<=26'd11304366; ROM3[3777]<=26'd9754188; ROM4[3777]<=26'd23471530;
ROM1[3778]<=26'd1987556; ROM2[3778]<=26'd11303598; ROM3[3778]<=26'd9758807; ROM4[3778]<=26'd23474112;
ROM1[3779]<=26'd1976553; ROM2[3779]<=26'd11296667; ROM3[3779]<=26'd9756044; ROM4[3779]<=26'd23469595;
ROM1[3780]<=26'd1979677; ROM2[3780]<=26'd11297116; ROM3[3780]<=26'd9756601; ROM4[3780]<=26'd23471733;
ROM1[3781]<=26'd1992218; ROM2[3781]<=26'd11300250; ROM3[3781]<=26'd9754933; ROM4[3781]<=26'd23474297;
ROM1[3782]<=26'd2003066; ROM2[3782]<=26'd11298753; ROM3[3782]<=26'd9746521; ROM4[3782]<=26'd23471389;
ROM1[3783]<=26'd2006831; ROM2[3783]<=26'd11299039; ROM3[3783]<=26'd9744092; ROM4[3783]<=26'd23472213;
ROM1[3784]<=26'd2001008; ROM2[3784]<=26'd11299484; ROM3[3784]<=26'd9747268; ROM4[3784]<=26'd23474005;
ROM1[3785]<=26'd1991998; ROM2[3785]<=26'd11298318; ROM3[3785]<=26'd9748383; ROM4[3785]<=26'd23473133;
ROM1[3786]<=26'd1987060; ROM2[3786]<=26'd11297258; ROM3[3786]<=26'd9748282; ROM4[3786]<=26'd23471170;
ROM1[3787]<=26'd1984166; ROM2[3787]<=26'd11295867; ROM3[3787]<=26'd9750212; ROM4[3787]<=26'd23470877;
ROM1[3788]<=26'd1986503; ROM2[3788]<=26'd11296606; ROM3[3788]<=26'd9753083; ROM4[3788]<=26'd23471908;
ROM1[3789]<=26'd1993185; ROM2[3789]<=26'd11299794; ROM3[3789]<=26'd9756692; ROM4[3789]<=26'd23474532;
ROM1[3790]<=26'd2002479; ROM2[3790]<=26'd11298391; ROM3[3790]<=26'd9753035; ROM4[3790]<=26'd23473688;
ROM1[3791]<=26'd2013379; ROM2[3791]<=26'd11302889; ROM3[3791]<=26'd9750612; ROM4[3791]<=26'd23475465;
ROM1[3792]<=26'd2014792; ROM2[3792]<=26'd11310458; ROM3[3792]<=26'd9755767; ROM4[3792]<=26'd23480971;
ROM1[3793]<=26'd2002411; ROM2[3793]<=26'd11303358; ROM3[3793]<=26'd9753692; ROM4[3793]<=26'd23475008;
ROM1[3794]<=26'd1985236; ROM2[3794]<=26'd11291576; ROM3[3794]<=26'd9747033; ROM4[3794]<=26'd23464688;
ROM1[3795]<=26'd1977495; ROM2[3795]<=26'd11289369; ROM3[3795]<=26'd9748987; ROM4[3795]<=26'd23463001;
ROM1[3796]<=26'd1970586; ROM2[3796]<=26'd11285543; ROM3[3796]<=26'd9747149; ROM4[3796]<=26'd23459133;
ROM1[3797]<=26'd1970983; ROM2[3797]<=26'd11283264; ROM3[3797]<=26'd9742154; ROM4[3797]<=26'd23455900;
ROM1[3798]<=26'd1985473; ROM2[3798]<=26'd11291335; ROM3[3798]<=26'd9742519; ROM4[3798]<=26'd23459929;
ROM1[3799]<=26'd1996668; ROM2[3799]<=26'd11292793; ROM3[3799]<=26'd9736386; ROM4[3799]<=26'd23460070;
ROM1[3800]<=26'd1995136; ROM2[3800]<=26'd11288996; ROM3[3800]<=26'd9734382; ROM4[3800]<=26'd23458082;
ROM1[3801]<=26'd1990545; ROM2[3801]<=26'd11290848; ROM3[3801]<=26'd9740168; ROM4[3801]<=26'd23461469;
ROM1[3802]<=26'd1986128; ROM2[3802]<=26'd11293997; ROM3[3802]<=26'd9746430; ROM4[3802]<=26'd23465638;
ROM1[3803]<=26'd1978469; ROM2[3803]<=26'd11291963; ROM3[3803]<=26'd9745220; ROM4[3803]<=26'd23463373;
ROM1[3804]<=26'd1968605; ROM2[3804]<=26'd11287988; ROM3[3804]<=26'd9742232; ROM4[3804]<=26'd23459504;
ROM1[3805]<=26'd1968016; ROM2[3805]<=26'd11287818; ROM3[3805]<=26'd9741356; ROM4[3805]<=26'd23459004;
ROM1[3806]<=26'd1974064; ROM2[3806]<=26'd11287129; ROM3[3806]<=26'd9736070; ROM4[3806]<=26'd23457208;
ROM1[3807]<=26'd1986058; ROM2[3807]<=26'd11289331; ROM3[3807]<=26'd9732255; ROM4[3807]<=26'd23457161;
ROM1[3808]<=26'd1993469; ROM2[3808]<=26'd11292105; ROM3[3808]<=26'd9733742; ROM4[3808]<=26'd23460427;
ROM1[3809]<=26'd1991810; ROM2[3809]<=26'd11294944; ROM3[3809]<=26'd9737740; ROM4[3809]<=26'd23462353;
ROM1[3810]<=26'd1990992; ROM2[3810]<=26'd11301885; ROM3[3810]<=26'd9748298; ROM4[3810]<=26'd23469557;
ROM1[3811]<=26'd1985547; ROM2[3811]<=26'd11300323; ROM3[3811]<=26'd9750494; ROM4[3811]<=26'd23470483;
ROM1[3812]<=26'd1969276; ROM2[3812]<=26'd11290782; ROM3[3812]<=26'd9741876; ROM4[3812]<=26'd23461419;
ROM1[3813]<=26'd1965928; ROM2[3813]<=26'd11288487; ROM3[3813]<=26'd9742846; ROM4[3813]<=26'd23461856;
ROM1[3814]<=26'd1974530; ROM2[3814]<=26'd11290558; ROM3[3814]<=26'd9743833; ROM4[3814]<=26'd23465336;
ROM1[3815]<=26'd1989171; ROM2[3815]<=26'd11291388; ROM3[3815]<=26'd9739983; ROM4[3815]<=26'd23465864;
ROM1[3816]<=26'd2003662; ROM2[3816]<=26'd11296602; ROM3[3816]<=26'd9742081; ROM4[3816]<=26'd23471339;
ROM1[3817]<=26'd2000142; ROM2[3817]<=26'd11297335; ROM3[3817]<=26'd9742217; ROM4[3817]<=26'd23471093;
ROM1[3818]<=26'd1991274; ROM2[3818]<=26'd11294225; ROM3[3818]<=26'd9741841; ROM4[3818]<=26'd23468957;
ROM1[3819]<=26'd1988103; ROM2[3819]<=26'd11296486; ROM3[3819]<=26'd9747731; ROM4[3819]<=26'd23471211;
ROM1[3820]<=26'd1984410; ROM2[3820]<=26'd11298327; ROM3[3820]<=26'd9751044; ROM4[3820]<=26'd23472343;
ROM1[3821]<=26'd1979289; ROM2[3821]<=26'd11296503; ROM3[3821]<=26'd9751290; ROM4[3821]<=26'd23469654;
ROM1[3822]<=26'd1978753; ROM2[3822]<=26'd11295359; ROM3[3822]<=26'd9747235; ROM4[3822]<=26'd23465544;
ROM1[3823]<=26'd1988195; ROM2[3823]<=26'd11297877; ROM3[3823]<=26'd9743678; ROM4[3823]<=26'd23466760;
ROM1[3824]<=26'd2002322; ROM2[3824]<=26'd11300590; ROM3[3824]<=26'd9741906; ROM4[3824]<=26'd23468265;
ROM1[3825]<=26'd1996758; ROM2[3825]<=26'd11295466; ROM3[3825]<=26'd9735651; ROM4[3825]<=26'd23463368;
ROM1[3826]<=26'd1989341; ROM2[3826]<=26'd11293814; ROM3[3826]<=26'd9737268; ROM4[3826]<=26'd23462971;
ROM1[3827]<=26'd1981570; ROM2[3827]<=26'd11292383; ROM3[3827]<=26'd9740093; ROM4[3827]<=26'd23462905;
ROM1[3828]<=26'd1974282; ROM2[3828]<=26'd11289910; ROM3[3828]<=26'd9742549; ROM4[3828]<=26'd23462624;
ROM1[3829]<=26'd1971715; ROM2[3829]<=26'd11291319; ROM3[3829]<=26'd9747717; ROM4[3829]<=26'd23465219;
ROM1[3830]<=26'd1972766; ROM2[3830]<=26'd11291034; ROM3[3830]<=26'd9747908; ROM4[3830]<=26'd23465660;
ROM1[3831]<=26'd1982306; ROM2[3831]<=26'd11290372; ROM3[3831]<=26'd9746244; ROM4[3831]<=26'd23464582;
ROM1[3832]<=26'd1995075; ROM2[3832]<=26'd11289933; ROM3[3832]<=26'd9739182; ROM4[3832]<=26'd23462059;
ROM1[3833]<=26'd2002430; ROM2[3833]<=26'd11291665; ROM3[3833]<=26'd9738306; ROM4[3833]<=26'd23465027;
ROM1[3834]<=26'd1995254; ROM2[3834]<=26'd11289440; ROM3[3834]<=26'd9742260; ROM4[3834]<=26'd23465907;
ROM1[3835]<=26'd1983293; ROM2[3835]<=26'd11284876; ROM3[3835]<=26'd9742581; ROM4[3835]<=26'd23463032;
ROM1[3836]<=26'd1983992; ROM2[3836]<=26'd11290216; ROM3[3836]<=26'd9749728; ROM4[3836]<=26'd23468208;
ROM1[3837]<=26'd1978579; ROM2[3837]<=26'd11290699; ROM3[3837]<=26'd9753294; ROM4[3837]<=26'd23469845;
ROM1[3838]<=26'd1970424; ROM2[3838]<=26'd11283276; ROM3[3838]<=26'd9747345; ROM4[3838]<=26'd23463790;
ROM1[3839]<=26'd1981026; ROM2[3839]<=26'd11289135; ROM3[3839]<=26'd9752057; ROM4[3839]<=26'd23468531;
ROM1[3840]<=26'd1991501; ROM2[3840]<=26'd11290169; ROM3[3840]<=26'd9748798; ROM4[3840]<=26'd23468352;
ROM1[3841]<=26'd1990959; ROM2[3841]<=26'd11282367; ROM3[3841]<=26'd9735344; ROM4[3841]<=26'd23458829;
ROM1[3842]<=26'd1991895; ROM2[3842]<=26'd11287405; ROM3[3842]<=26'd9739291; ROM4[3842]<=26'd23462677;
ROM1[3843]<=26'd1984657; ROM2[3843]<=26'd11287638; ROM3[3843]<=26'd9741955; ROM4[3843]<=26'd23463568;
ROM1[3844]<=26'd1974849; ROM2[3844]<=26'd11284593; ROM3[3844]<=26'd9741473; ROM4[3844]<=26'd23460797;
ROM1[3845]<=26'd1973454; ROM2[3845]<=26'd11288568; ROM3[3845]<=26'd9747094; ROM4[3845]<=26'd23465533;
ROM1[3846]<=26'd1970030; ROM2[3846]<=26'd11289103; ROM3[3846]<=26'd9750024; ROM4[3846]<=26'd23466914;
ROM1[3847]<=26'd1972310; ROM2[3847]<=26'd11290377; ROM3[3847]<=26'd9748518; ROM4[3847]<=26'd23465704;
ROM1[3848]<=26'd1984550; ROM2[3848]<=26'd11291995; ROM3[3848]<=26'd9744568; ROM4[3848]<=26'd23466575;
ROM1[3849]<=26'd2001397; ROM2[3849]<=26'd11296548; ROM3[3849]<=26'd9744990; ROM4[3849]<=26'd23470746;
ROM1[3850]<=26'd2004784; ROM2[3850]<=26'd11298346; ROM3[3850]<=26'd9744592; ROM4[3850]<=26'd23471683;
ROM1[3851]<=26'd1998214; ROM2[3851]<=26'd11296942; ROM3[3851]<=26'd9745752; ROM4[3851]<=26'd23470934;
ROM1[3852]<=26'd1989167; ROM2[3852]<=26'd11295941; ROM3[3852]<=26'd9748699; ROM4[3852]<=26'd23468531;
ROM1[3853]<=26'd1983162; ROM2[3853]<=26'd11295442; ROM3[3853]<=26'd9750272; ROM4[3853]<=26'd23466120;
ROM1[3854]<=26'd1975050; ROM2[3854]<=26'd11293047; ROM3[3854]<=26'd9750320; ROM4[3854]<=26'd23464250;
ROM1[3855]<=26'd1972426; ROM2[3855]<=26'd11290827; ROM3[3855]<=26'd9747952; ROM4[3855]<=26'd23463200;
ROM1[3856]<=26'd1983529; ROM2[3856]<=26'd11294046; ROM3[3856]<=26'd9746907; ROM4[3856]<=26'd23465709;
ROM1[3857]<=26'd1998934; ROM2[3857]<=26'd11296888; ROM3[3857]<=26'd9744300; ROM4[3857]<=26'd23468381;
ROM1[3858]<=26'd2003828; ROM2[3858]<=26'd11296961; ROM3[3858]<=26'd9741835; ROM4[3858]<=26'd23467233;
ROM1[3859]<=26'd1999169; ROM2[3859]<=26'd11296675; ROM3[3859]<=26'd9744250; ROM4[3859]<=26'd23467211;
ROM1[3860]<=26'd1992954; ROM2[3860]<=26'd11297373; ROM3[3860]<=26'd9749606; ROM4[3860]<=26'd23470889;
ROM1[3861]<=26'd1988592; ROM2[3861]<=26'd11296681; ROM3[3861]<=26'd9751935; ROM4[3861]<=26'd23471837;
ROM1[3862]<=26'd1983793; ROM2[3862]<=26'd11296285; ROM3[3862]<=26'd9755071; ROM4[3862]<=26'd23473130;
ROM1[3863]<=26'd1980383; ROM2[3863]<=26'd11294500; ROM3[3863]<=26'd9755508; ROM4[3863]<=26'd23472803;
ROM1[3864]<=26'd1981865; ROM2[3864]<=26'd11290826; ROM3[3864]<=26'd9751187; ROM4[3864]<=26'd23470368;
ROM1[3865]<=26'd1993790; ROM2[3865]<=26'd11292675; ROM3[3865]<=26'd9748615; ROM4[3865]<=26'd23471957;
ROM1[3866]<=26'd2013149; ROM2[3866]<=26'd11303742; ROM3[3866]<=26'd9753885; ROM4[3866]<=26'd23480813;
ROM1[3867]<=26'd2012486; ROM2[3867]<=26'd11303549; ROM3[3867]<=26'd9754780; ROM4[3867]<=26'd23481608;
ROM1[3868]<=26'd1995652; ROM2[3868]<=26'd11290714; ROM3[3868]<=26'd9746764; ROM4[3868]<=26'd23470280;
ROM1[3869]<=26'd1986575; ROM2[3869]<=26'd11287704; ROM3[3869]<=26'd9746963; ROM4[3869]<=26'd23466603;
ROM1[3870]<=26'd1978407; ROM2[3870]<=26'd11284409; ROM3[3870]<=26'd9747209; ROM4[3870]<=26'd23464451;
ROM1[3871]<=26'd1971940; ROM2[3871]<=26'd11281487; ROM3[3871]<=26'd9746305; ROM4[3871]<=26'd23462007;
ROM1[3872]<=26'd1981366; ROM2[3872]<=26'd11287697; ROM3[3872]<=26'd9750576; ROM4[3872]<=26'd23467408;
ROM1[3873]<=26'd1997835; ROM2[3873]<=26'd11294483; ROM3[3873]<=26'd9753412; ROM4[3873]<=26'd23472981;
ROM1[3874]<=26'd2010634; ROM2[3874]<=26'd11296588; ROM3[3874]<=26'd9748658; ROM4[3874]<=26'd23471754;
ROM1[3875]<=26'd2012259; ROM2[3875]<=26'd11297263; ROM3[3875]<=26'd9748174; ROM4[3875]<=26'd23471632;
ROM1[3876]<=26'd2004262; ROM2[3876]<=26'd11296961; ROM3[3876]<=26'd9753258; ROM4[3876]<=26'd23473323;
ROM1[3877]<=26'd1993250; ROM2[3877]<=26'd11291359; ROM3[3877]<=26'd9753871; ROM4[3877]<=26'd23470253;
ROM1[3878]<=26'd1986179; ROM2[3878]<=26'd11289779; ROM3[3878]<=26'd9755460; ROM4[3878]<=26'd23469634;
ROM1[3879]<=26'd1984665; ROM2[3879]<=26'd11294333; ROM3[3879]<=26'd9759911; ROM4[3879]<=26'd23473216;
ROM1[3880]<=26'd1992049; ROM2[3880]<=26'd11302586; ROM3[3880]<=26'd9762511; ROM4[3880]<=26'd23479430;
ROM1[3881]<=26'd1999174; ROM2[3881]<=26'd11303964; ROM3[3881]<=26'd9756725; ROM4[3881]<=26'd23479210;
ROM1[3882]<=26'd2007189; ROM2[3882]<=26'd11298546; ROM3[3882]<=26'd9746768; ROM4[3882]<=26'd23474373;
ROM1[3883]<=26'd2012000; ROM2[3883]<=26'd11299136; ROM3[3883]<=26'd9744633; ROM4[3883]<=26'd23474376;
ROM1[3884]<=26'd2009807; ROM2[3884]<=26'd11301996; ROM3[3884]<=26'd9749559; ROM4[3884]<=26'd23477409;
ROM1[3885]<=26'd1999076; ROM2[3885]<=26'd11296387; ROM3[3885]<=26'd9750952; ROM4[3885]<=26'd23474520;
ROM1[3886]<=26'd1992191; ROM2[3886]<=26'd11295732; ROM3[3886]<=26'd9753763; ROM4[3886]<=26'd23475900;
ROM1[3887]<=26'd1988817; ROM2[3887]<=26'd11297966; ROM3[3887]<=26'd9760543; ROM4[3887]<=26'd23481576;
ROM1[3888]<=26'd1992200; ROM2[3888]<=26'd11302096; ROM3[3888]<=26'd9766760; ROM4[3888]<=26'd23486830;
ROM1[3889]<=26'd1997637; ROM2[3889]<=26'd11303200; ROM3[3889]<=26'd9764630; ROM4[3889]<=26'd23486650;
ROM1[3890]<=26'd2003163; ROM2[3890]<=26'd11296937; ROM3[3890]<=26'd9753838; ROM4[3890]<=26'd23478040;
ROM1[3891]<=26'd2005688; ROM2[3891]<=26'd11291989; ROM3[3891]<=26'd9743256; ROM4[3891]<=26'd23470943;
ROM1[3892]<=26'd1999349; ROM2[3892]<=26'd11290024; ROM3[3892]<=26'd9742559; ROM4[3892]<=26'd23468907;
ROM1[3893]<=26'd1998622; ROM2[3893]<=26'd11297297; ROM3[3893]<=26'd9752261; ROM4[3893]<=26'd23476058;
ROM1[3894]<=26'd1996680; ROM2[3894]<=26'd11301256; ROM3[3894]<=26'd9760669; ROM4[3894]<=26'd23481485;
ROM1[3895]<=26'd1988178; ROM2[3895]<=26'd11299484; ROM3[3895]<=26'd9762850; ROM4[3895]<=26'd23479833;
ROM1[3896]<=26'd1977236; ROM2[3896]<=26'd11292951; ROM3[3896]<=26'd9759107; ROM4[3896]<=26'd23474464;
ROM1[3897]<=26'd1975516; ROM2[3897]<=26'd11286709; ROM3[3897]<=26'd9753639; ROM4[3897]<=26'd23470365;
ROM1[3898]<=26'd1982466; ROM2[3898]<=26'd11284704; ROM3[3898]<=26'd9747555; ROM4[3898]<=26'd23467980;
ROM1[3899]<=26'd1996934; ROM2[3899]<=26'd11288150; ROM3[3899]<=26'd9745095; ROM4[3899]<=26'd23470995;
ROM1[3900]<=26'd2002704; ROM2[3900]<=26'd11293206; ROM3[3900]<=26'd9746042; ROM4[3900]<=26'd23473904;
ROM1[3901]<=26'd1995049; ROM2[3901]<=26'd11293915; ROM3[3901]<=26'd9743553; ROM4[3901]<=26'd23469722;
ROM1[3902]<=26'd1988198; ROM2[3902]<=26'd11293372; ROM3[3902]<=26'd9741432; ROM4[3902]<=26'd23467157;
ROM1[3903]<=26'd1985947; ROM2[3903]<=26'd11294179; ROM3[3903]<=26'd9744492; ROM4[3903]<=26'd23470402;
ROM1[3904]<=26'd1979371; ROM2[3904]<=26'd11295990; ROM3[3904]<=26'd9747843; ROM4[3904]<=26'd23473778;
ROM1[3905]<=26'd1981572; ROM2[3905]<=26'd11299437; ROM3[3905]<=26'd9751665; ROM4[3905]<=26'd23476313;
ROM1[3906]<=26'd2000852; ROM2[3906]<=26'd11311257; ROM3[3906]<=26'd9759022; ROM4[3906]<=26'd23485232;
ROM1[3907]<=26'd2018396; ROM2[3907]<=26'd11316043; ROM3[3907]<=26'd9757609; ROM4[3907]<=26'd23488198;
ROM1[3908]<=26'd2015585; ROM2[3908]<=26'd11307435; ROM3[3908]<=26'd9747717; ROM4[3908]<=26'd23477784;
ROM1[3909]<=26'd2010617; ROM2[3909]<=26'd11307826; ROM3[3909]<=26'd9750666; ROM4[3909]<=26'd23478211;
ROM1[3910]<=26'd2003327; ROM2[3910]<=26'd11306738; ROM3[3910]<=26'd9754644; ROM4[3910]<=26'd23480458;
ROM1[3911]<=26'd1995536; ROM2[3911]<=26'd11304977; ROM3[3911]<=26'd9753462; ROM4[3911]<=26'd23476103;
ROM1[3912]<=26'd1994119; ROM2[3912]<=26'd11307074; ROM3[3912]<=26'd9758559; ROM4[3912]<=26'd23478289;
ROM1[3913]<=26'd1991532; ROM2[3913]<=26'd11306177; ROM3[3913]<=26'd9761741; ROM4[3913]<=26'd23480852;
ROM1[3914]<=26'd1993364; ROM2[3914]<=26'd11304659; ROM3[3914]<=26'd9758088; ROM4[3914]<=26'd23479613;
ROM1[3915]<=26'd2003525; ROM2[3915]<=26'd11304431; ROM3[3915]<=26'd9752813; ROM4[3915]<=26'd23478529;
ROM1[3916]<=26'd2013170; ROM2[3916]<=26'd11306449; ROM3[3916]<=26'd9751001; ROM4[3916]<=26'd23479415;
ROM1[3917]<=26'd2010568; ROM2[3917]<=26'd11306036; ROM3[3917]<=26'd9751559; ROM4[3917]<=26'd23480607;
ROM1[3918]<=26'd2002881; ROM2[3918]<=26'd11304523; ROM3[3918]<=26'd9755594; ROM4[3918]<=26'd23482824;
ROM1[3919]<=26'd1996852; ROM2[3919]<=26'd11303988; ROM3[3919]<=26'd9760626; ROM4[3919]<=26'd23483829;
ROM1[3920]<=26'd1991449; ROM2[3920]<=26'd11303771; ROM3[3920]<=26'd9763403; ROM4[3920]<=26'd23484272;
ROM1[3921]<=26'd1989744; ROM2[3921]<=26'd11305353; ROM3[3921]<=26'd9768029; ROM4[3921]<=26'd23485470;
ROM1[3922]<=26'd1997524; ROM2[3922]<=26'd11310979; ROM3[3922]<=26'd9770051; ROM4[3922]<=26'd23486677;
ROM1[3923]<=26'd2010928; ROM2[3923]<=26'd11315441; ROM3[3923]<=26'd9768418; ROM4[3923]<=26'd23489355;
ROM1[3924]<=26'd2024718; ROM2[3924]<=26'd11319672; ROM3[3924]<=26'd9768253; ROM4[3924]<=26'd23492598;
ROM1[3925]<=26'd2017517; ROM2[3925]<=26'd11312975; ROM3[3925]<=26'd9758907; ROM4[3925]<=26'd23485171;
ROM1[3926]<=26'd2006998; ROM2[3926]<=26'd11309058; ROM3[3926]<=26'd9758674; ROM4[3926]<=26'd23481363;
ROM1[3927]<=26'd2003262; ROM2[3927]<=26'd11312548; ROM3[3927]<=26'd9764540; ROM4[3927]<=26'd23484386;
ROM1[3928]<=26'd1999068; ROM2[3928]<=26'd11312024; ROM3[3928]<=26'd9764666; ROM4[3928]<=26'd23485259;
ROM1[3929]<=26'd1990910; ROM2[3929]<=26'd11307999; ROM3[3929]<=26'd9765010; ROM4[3929]<=26'd23483333;
ROM1[3930]<=26'd1988356; ROM2[3930]<=26'd11307545; ROM3[3930]<=26'd9763579; ROM4[3930]<=26'd23483051;
ROM1[3931]<=26'd1991605; ROM2[3931]<=26'd11305099; ROM3[3931]<=26'd9757503; ROM4[3931]<=26'd23481544;
ROM1[3932]<=26'd2001953; ROM2[3932]<=26'd11303263; ROM3[3932]<=26'd9749167; ROM4[3932]<=26'd23478584;
ROM1[3933]<=26'd2011366; ROM2[3933]<=26'd11308039; ROM3[3933]<=26'd9749283; ROM4[3933]<=26'd23482420;
ROM1[3934]<=26'd2005964; ROM2[3934]<=26'd11307042; ROM3[3934]<=26'd9751845; ROM4[3934]<=26'd23482823;
ROM1[3935]<=26'd1998270; ROM2[3935]<=26'd11303299; ROM3[3935]<=26'd9754613; ROM4[3935]<=26'd23481582;
ROM1[3936]<=26'd1992975; ROM2[3936]<=26'd11303351; ROM3[3936]<=26'd9756423; ROM4[3936]<=26'd23481319;
ROM1[3937]<=26'd1990082; ROM2[3937]<=26'd11305916; ROM3[3937]<=26'd9762506; ROM4[3937]<=26'd23483061;
ROM1[3938]<=26'd1987688; ROM2[3938]<=26'd11305470; ROM3[3938]<=26'd9764396; ROM4[3938]<=26'd23483607;
ROM1[3939]<=26'd1988504; ROM2[3939]<=26'd11303920; ROM3[3939]<=26'd9759572; ROM4[3939]<=26'd23480399;
ROM1[3940]<=26'd1998874; ROM2[3940]<=26'd11303200; ROM3[3940]<=26'd9755048; ROM4[3940]<=26'd23478554;
ROM1[3941]<=26'd2009909; ROM2[3941]<=26'd11306232; ROM3[3941]<=26'd9753704; ROM4[3941]<=26'd23480790;
ROM1[3942]<=26'd2012067; ROM2[3942]<=26'd11309995; ROM3[3942]<=26'd9759261; ROM4[3942]<=26'd23485187;
ROM1[3943]<=26'd2003119; ROM2[3943]<=26'd11308573; ROM3[3943]<=26'd9760981; ROM4[3943]<=26'd23483086;
ROM1[3944]<=26'd1992603; ROM2[3944]<=26'd11304191; ROM3[3944]<=26'd9761935; ROM4[3944]<=26'd23478560;
ROM1[3945]<=26'd1986562; ROM2[3945]<=26'd11301807; ROM3[3945]<=26'd9762695; ROM4[3945]<=26'd23477357;
ROM1[3946]<=26'd1977842; ROM2[3946]<=26'd11297162; ROM3[3946]<=26'd9758635; ROM4[3946]<=26'd23472833;
ROM1[3947]<=26'd1985964; ROM2[3947]<=26'd11302573; ROM3[3947]<=26'd9762352; ROM4[3947]<=26'd23477404;
ROM1[3948]<=26'd2003456; ROM2[3948]<=26'd11309777; ROM3[3948]<=26'd9764416; ROM4[3948]<=26'd23484090;
ROM1[3949]<=26'd2009531; ROM2[3949]<=26'd11304504; ROM3[3949]<=26'd9753869; ROM4[3949]<=26'd23479664;
ROM1[3950]<=26'd2007496; ROM2[3950]<=26'd11302123; ROM3[3950]<=26'd9750108; ROM4[3950]<=26'd23476163;
ROM1[3951]<=26'd1997561; ROM2[3951]<=26'd11299790; ROM3[3951]<=26'd9752240; ROM4[3951]<=26'd23474126;
ROM1[3952]<=26'd1989999; ROM2[3952]<=26'd11297102; ROM3[3952]<=26'd9753596; ROM4[3952]<=26'd23473902;
ROM1[3953]<=26'd1989065; ROM2[3953]<=26'd11300463; ROM3[3953]<=26'd9759067; ROM4[3953]<=26'd23479145;
ROM1[3954]<=26'd1986696; ROM2[3954]<=26'd11303078; ROM3[3954]<=26'd9763679; ROM4[3954]<=26'd23482766;
ROM1[3955]<=26'd1989734; ROM2[3955]<=26'd11304713; ROM3[3955]<=26'd9765367; ROM4[3955]<=26'd23485429;
ROM1[3956]<=26'd1993503; ROM2[3956]<=26'd11302261; ROM3[3956]<=26'd9758386; ROM4[3956]<=26'd23482637;
ROM1[3957]<=26'd1999850; ROM2[3957]<=26'd11297948; ROM3[3957]<=26'd9747504; ROM4[3957]<=26'd23475615;
ROM1[3958]<=26'd2003638; ROM2[3958]<=26'd11297138; ROM3[3958]<=26'd9744930; ROM4[3958]<=26'd23475796;
ROM1[3959]<=26'd2001537; ROM2[3959]<=26'd11297246; ROM3[3959]<=26'd9747284; ROM4[3959]<=26'd23478233;
ROM1[3960]<=26'd2001465; ROM2[3960]<=26'd11302658; ROM3[3960]<=26'd9757113; ROM4[3960]<=26'd23483136;
ROM1[3961]<=26'd1999174; ROM2[3961]<=26'd11305430; ROM3[3961]<=26'd9763487; ROM4[3961]<=26'd23486824;
ROM1[3962]<=26'd1988643; ROM2[3962]<=26'd11300376; ROM3[3962]<=26'd9760648; ROM4[3962]<=26'd23483253;
ROM1[3963]<=26'd1981543; ROM2[3963]<=26'd11295211; ROM3[3963]<=26'd9757304; ROM4[3963]<=26'd23478099;
ROM1[3964]<=26'd1985725; ROM2[3964]<=26'd11295371; ROM3[3964]<=26'd9754636; ROM4[3964]<=26'd23477715;
ROM1[3965]<=26'd2000578; ROM2[3965]<=26'd11301457; ROM3[3965]<=26'd9750473; ROM4[3965]<=26'd23480840;
ROM1[3966]<=26'd2009429; ROM2[3966]<=26'd11301190; ROM3[3966]<=26'd9744290; ROM4[3966]<=26'd23478742;
ROM1[3967]<=26'd2003475; ROM2[3967]<=26'd11297908; ROM3[3967]<=26'd9741409; ROM4[3967]<=26'd23474876;
ROM1[3968]<=26'd1992843; ROM2[3968]<=26'd11295737; ROM3[3968]<=26'd9743901; ROM4[3968]<=26'd23474253;
ROM1[3969]<=26'd1990818; ROM2[3969]<=26'd11298563; ROM3[3969]<=26'd9753217; ROM4[3969]<=26'd23479543;
ROM1[3970]<=26'd1995336; ROM2[3970]<=26'd11307292; ROM3[3970]<=26'd9765243; ROM4[3970]<=26'd23489496;
ROM1[3971]<=26'd1997623; ROM2[3971]<=26'd11311614; ROM3[3971]<=26'd9772596; ROM4[3971]<=26'd23493806;
ROM1[3972]<=26'd2000137; ROM2[3972]<=26'd11310577; ROM3[3972]<=26'd9770462; ROM4[3972]<=26'd23490884;
ROM1[3973]<=26'd2007083; ROM2[3973]<=26'd11308492; ROM3[3973]<=26'd9765530; ROM4[3973]<=26'd23487654;
ROM1[3974]<=26'd2013919; ROM2[3974]<=26'd11306883; ROM3[3974]<=26'd9761140; ROM4[3974]<=26'd23484515;
ROM1[3975]<=26'd2011868; ROM2[3975]<=26'd11306645; ROM3[3975]<=26'd9758826; ROM4[3975]<=26'd23483689;
ROM1[3976]<=26'd2010266; ROM2[3976]<=26'd11308347; ROM3[3976]<=26'd9764473; ROM4[3976]<=26'd23489067;
ROM1[3977]<=26'd2001380; ROM2[3977]<=26'd11304627; ROM3[3977]<=26'd9765876; ROM4[3977]<=26'd23485965;
ROM1[3978]<=26'd1992757; ROM2[3978]<=26'd11300454; ROM3[3978]<=26'd9765152; ROM4[3978]<=26'd23481752;
ROM1[3979]<=26'd1987115; ROM2[3979]<=26'd11298207; ROM3[3979]<=26'd9767988; ROM4[3979]<=26'd23481094;
ROM1[3980]<=26'd1990529; ROM2[3980]<=26'd11302710; ROM3[3980]<=26'd9770631; ROM4[3980]<=26'd23484413;
ROM1[3981]<=26'd2007562; ROM2[3981]<=26'd11314402; ROM3[3981]<=26'd9775776; ROM4[3981]<=26'd23492621;
ROM1[3982]<=26'd2018572; ROM2[3982]<=26'd11313590; ROM3[3982]<=26'd9768319; ROM4[3982]<=26'd23490075;
ROM1[3983]<=26'd2016317; ROM2[3983]<=26'd11308428; ROM3[3983]<=26'd9757014; ROM4[3983]<=26'd23483580;
ROM1[3984]<=26'd2010778; ROM2[3984]<=26'd11309840; ROM3[3984]<=26'd9758002; ROM4[3984]<=26'd23482712;
ROM1[3985]<=26'd2000873; ROM2[3985]<=26'd11307192; ROM3[3985]<=26'd9759600; ROM4[3985]<=26'd23480880;
ROM1[3986]<=26'd1993047; ROM2[3986]<=26'd11304648; ROM3[3986]<=26'd9759599; ROM4[3986]<=26'd23480001;
ROM1[3987]<=26'd1985752; ROM2[3987]<=26'd11302122; ROM3[3987]<=26'd9760279; ROM4[3987]<=26'd23478190;
ROM1[3988]<=26'd1980289; ROM2[3988]<=26'd11298561; ROM3[3988]<=26'd9758315; ROM4[3988]<=26'd23476235;
ROM1[3989]<=26'd1984877; ROM2[3989]<=26'd11297337; ROM3[3989]<=26'd9753263; ROM4[3989]<=26'd23474174;
ROM1[3990]<=26'd2000523; ROM2[3990]<=26'd11302954; ROM3[3990]<=26'd9751628; ROM4[3990]<=26'd23475771;
ROM1[3991]<=26'd2014124; ROM2[3991]<=26'd11308577; ROM3[3991]<=26'd9751658; ROM4[3991]<=26'd23481061;
ROM1[3992]<=26'd2007251; ROM2[3992]<=26'd11305328; ROM3[3992]<=26'd9749594; ROM4[3992]<=26'd23479405;
ROM1[3993]<=26'd2000152; ROM2[3993]<=26'd11306294; ROM3[3993]<=26'd9753269; ROM4[3993]<=26'd23480894;
ROM1[3994]<=26'd2000854; ROM2[3994]<=26'd11311825; ROM3[3994]<=26'd9761350; ROM4[3994]<=26'd23486907;
ROM1[3995]<=26'd1997664; ROM2[3995]<=26'd11314064; ROM3[3995]<=26'd9766307; ROM4[3995]<=26'd23489592;
ROM1[3996]<=26'd1992328; ROM2[3996]<=26'd11311984; ROM3[3996]<=26'd9765872; ROM4[3996]<=26'd23488017;
ROM1[3997]<=26'd1989499; ROM2[3997]<=26'd11305800; ROM3[3997]<=26'd9760154; ROM4[3997]<=26'd23480573;
ROM1[3998]<=26'd1992287; ROM2[3998]<=26'd11298958; ROM3[3998]<=26'd9749412; ROM4[3998]<=26'd23472618;
ROM1[3999]<=26'd2002362; ROM2[3999]<=26'd11298970; ROM3[3999]<=26'd9744105; ROM4[3999]<=26'd23470867;
ROM1[4000]<=26'd2001309; ROM2[4000]<=26'd11297053; ROM3[4000]<=26'd9742601; ROM4[4000]<=26'd23468218;
ROM1[4001]<=26'd1996374; ROM2[4001]<=26'd11295314; ROM3[4001]<=26'd9744646; ROM4[4001]<=26'd23470834;
ROM1[4002]<=26'd1991856; ROM2[4002]<=26'd11296809; ROM3[4002]<=26'd9751128; ROM4[4002]<=26'd23473625;
ROM1[4003]<=26'd1983411; ROM2[4003]<=26'd11293064; ROM3[4003]<=26'd9751309; ROM4[4003]<=26'd23471675;
ROM1[4004]<=26'd1976005; ROM2[4004]<=26'd11290125; ROM3[4004]<=26'd9752445; ROM4[4004]<=26'd23472005;
ROM1[4005]<=26'd1978075; ROM2[4005]<=26'd11293882; ROM3[4005]<=26'd9755998; ROM4[4005]<=26'd23474213;
ROM1[4006]<=26'd1989991; ROM2[4006]<=26'd11297028; ROM3[4006]<=26'd9755651; ROM4[4006]<=26'd23477459;
ROM1[4007]<=26'd2003540; ROM2[4007]<=26'd11296402; ROM3[4007]<=26'd9750238; ROM4[4007]<=26'd23477812;
ROM1[4008]<=26'd2008778; ROM2[4008]<=26'd11298752; ROM3[4008]<=26'd9748252; ROM4[4008]<=26'd23477943;
ROM1[4009]<=26'd2003100; ROM2[4009]<=26'd11297786; ROM3[4009]<=26'd9748951; ROM4[4009]<=26'd23477139;
ROM1[4010]<=26'd1991837; ROM2[4010]<=26'd11293884; ROM3[4010]<=26'd9748654; ROM4[4010]<=26'd23475168;
ROM1[4011]<=26'd1986203; ROM2[4011]<=26'd11295472; ROM3[4011]<=26'd9753162; ROM4[4011]<=26'd23475973;
ROM1[4012]<=26'd1983915; ROM2[4012]<=26'd11295886; ROM3[4012]<=26'd9757454; ROM4[4012]<=26'd23476321;
ROM1[4013]<=26'd1981123; ROM2[4013]<=26'd11294837; ROM3[4013]<=26'd9756719; ROM4[4013]<=26'd23475049;
ROM1[4014]<=26'd1990308; ROM2[4014]<=26'd11299380; ROM3[4014]<=26'd9759788; ROM4[4014]<=26'd23478771;
ROM1[4015]<=26'd2012504; ROM2[4015]<=26'd11310939; ROM3[4015]<=26'd9765955; ROM4[4015]<=26'd23490122;
ROM1[4016]<=26'd2020049; ROM2[4016]<=26'd11311889; ROM3[4016]<=26'd9761743; ROM4[4016]<=26'd23490536;
ROM1[4017]<=26'd2008966; ROM2[4017]<=26'd11303091; ROM3[4017]<=26'd9754680; ROM4[4017]<=26'd23482992;
ROM1[4018]<=26'd1994371; ROM2[4018]<=26'd11297980; ROM3[4018]<=26'd9751307; ROM4[4018]<=26'd23478035;
ROM1[4019]<=26'd1984254; ROM2[4019]<=26'd11295738; ROM3[4019]<=26'd9751191; ROM4[4019]<=26'd23474161;
ROM1[4020]<=26'd1981289; ROM2[4020]<=26'd11296386; ROM3[4020]<=26'd9753931; ROM4[4020]<=26'd23474270;
ROM1[4021]<=26'd1978572; ROM2[4021]<=26'd11297943; ROM3[4021]<=26'd9755999; ROM4[4021]<=26'd23474571;
ROM1[4022]<=26'd1981657; ROM2[4022]<=26'd11298824; ROM3[4022]<=26'd9755987; ROM4[4022]<=26'd23473285;
ROM1[4023]<=26'd1992693; ROM2[4023]<=26'd11298262; ROM3[4023]<=26'd9751625; ROM4[4023]<=26'd23472915;
ROM1[4024]<=26'd2001433; ROM2[4024]<=26'd11297329; ROM3[4024]<=26'd9744085; ROM4[4024]<=26'd23470371;
ROM1[4025]<=26'd2001777; ROM2[4025]<=26'd11297027; ROM3[4025]<=26'd9743256; ROM4[4025]<=26'd23469153;
ROM1[4026]<=26'd1997901; ROM2[4026]<=26'd11297654; ROM3[4026]<=26'd9745551; ROM4[4026]<=26'd23472264;
ROM1[4027]<=26'd1994101; ROM2[4027]<=26'd11301424; ROM3[4027]<=26'd9753234; ROM4[4027]<=26'd23475861;
ROM1[4028]<=26'd1988325; ROM2[4028]<=26'd11300620; ROM3[4028]<=26'd9756662; ROM4[4028]<=26'd23476021;
ROM1[4029]<=26'd1976599; ROM2[4029]<=26'd11294216; ROM3[4029]<=26'd9753576; ROM4[4029]<=26'd23471658;
ROM1[4030]<=26'd1977321; ROM2[4030]<=26'd11296595; ROM3[4030]<=26'd9751572; ROM4[4030]<=26'd23471768;
ROM1[4031]<=26'd1986194; ROM2[4031]<=26'd11296003; ROM3[4031]<=26'd9744640; ROM4[4031]<=26'd23469818;
ROM1[4032]<=26'd2006097; ROM2[4032]<=26'd11303137; ROM3[4032]<=26'd9747957; ROM4[4032]<=26'd23474957;
ROM1[4033]<=26'd2011547; ROM2[4033]<=26'd11305355; ROM3[4033]<=26'd9749004; ROM4[4033]<=26'd23477619;
ROM1[4034]<=26'd1993274; ROM2[4034]<=26'd11291754; ROM3[4034]<=26'd9742325; ROM4[4034]<=26'd23467045;
ROM1[4035]<=26'd1980996; ROM2[4035]<=26'd11286511; ROM3[4035]<=26'd9743764; ROM4[4035]<=26'd23463612;
ROM1[4036]<=26'd1973631; ROM2[4036]<=26'd11284080; ROM3[4036]<=26'd9744922; ROM4[4036]<=26'd23463102;
ROM1[4037]<=26'd1971298; ROM2[4037]<=26'd11286068; ROM3[4037]<=26'd9751338; ROM4[4037]<=26'd23466712;
ROM1[4038]<=26'd1977255; ROM2[4038]<=26'd11293205; ROM3[4038]<=26'd9760683; ROM4[4038]<=26'd23473870;
ROM1[4039]<=26'd1980178; ROM2[4039]<=26'd11290767; ROM3[4039]<=26'd9756739; ROM4[4039]<=26'd23470805;
ROM1[4040]<=26'd1988073; ROM2[4040]<=26'd11287726; ROM3[4040]<=26'd9746770; ROM4[4040]<=26'd23465674;
ROM1[4041]<=26'd2000923; ROM2[4041]<=26'd11291358; ROM3[4041]<=26'd9744504; ROM4[4041]<=26'd23467448;
ROM1[4042]<=26'd2001954; ROM2[4042]<=26'd11293217; ROM3[4042]<=26'd9746529; ROM4[4042]<=26'd23469051;
ROM1[4043]<=26'd1996107; ROM2[4043]<=26'd11294378; ROM3[4043]<=26'd9751088; ROM4[4043]<=26'd23470330;
ROM1[4044]<=26'd1991283; ROM2[4044]<=26'd11294840; ROM3[4044]<=26'd9757184; ROM4[4044]<=26'd23472121;
ROM1[4045]<=26'd1986770; ROM2[4045]<=26'd11295183; ROM3[4045]<=26'd9760995; ROM4[4045]<=26'd23473021;
ROM1[4046]<=26'd1981144; ROM2[4046]<=26'd11294165; ROM3[4046]<=26'd9761823; ROM4[4046]<=26'd23472459;
ROM1[4047]<=26'd1985720; ROM2[4047]<=26'd11296997; ROM3[4047]<=26'd9762296; ROM4[4047]<=26'd23475400;
ROM1[4048]<=26'd1994563; ROM2[4048]<=26'd11297195; ROM3[4048]<=26'd9755848; ROM4[4048]<=26'd23473651;
ROM1[4049]<=26'd2003026; ROM2[4049]<=26'd11296407; ROM3[4049]<=26'd9746200; ROM4[4049]<=26'd23471550;
ROM1[4050]<=26'd2007987; ROM2[4050]<=26'd11301308; ROM3[4050]<=26'd9748777; ROM4[4050]<=26'd23476341;
ROM1[4051]<=26'd2002013; ROM2[4051]<=26'd11301492; ROM3[4051]<=26'd9750938; ROM4[4051]<=26'd23475672;
ROM1[4052]<=26'd1991487; ROM2[4052]<=26'd11296512; ROM3[4052]<=26'd9748790; ROM4[4052]<=26'd23473602;
ROM1[4053]<=26'd1987948; ROM2[4053]<=26'd11295984; ROM3[4053]<=26'd9752354; ROM4[4053]<=26'd23474186;
ROM1[4054]<=26'd1983569; ROM2[4054]<=26'd11296611; ROM3[4054]<=26'd9756566; ROM4[4054]<=26'd23474680;
ROM1[4055]<=26'd1980256; ROM2[4055]<=26'd11293383; ROM3[4055]<=26'd9752890; ROM4[4055]<=26'd23471745;
ROM1[4056]<=26'd1989895; ROM2[4056]<=26'd11296874; ROM3[4056]<=26'd9751092; ROM4[4056]<=26'd23472914;
ROM1[4057]<=26'd2003764; ROM2[4057]<=26'd11300317; ROM3[4057]<=26'd9748548; ROM4[4057]<=26'd23475388;
ROM1[4058]<=26'd2004696; ROM2[4058]<=26'd11298048; ROM3[4058]<=26'd9744466; ROM4[4058]<=26'd23471661;
ROM1[4059]<=26'd1997906; ROM2[4059]<=26'd11295976; ROM3[4059]<=26'd9747237; ROM4[4059]<=26'd23471675;
ROM1[4060]<=26'd1991076; ROM2[4060]<=26'd11295591; ROM3[4060]<=26'd9752157; ROM4[4060]<=26'd23473237;
ROM1[4061]<=26'd1985369; ROM2[4061]<=26'd11295569; ROM3[4061]<=26'd9754735; ROM4[4061]<=26'd23472971;
ROM1[4062]<=26'd1976947; ROM2[4062]<=26'd11291410; ROM3[4062]<=26'd9753007; ROM4[4062]<=26'd23470261;
ROM1[4063]<=26'd1972483; ROM2[4063]<=26'd11288327; ROM3[4063]<=26'd9751058; ROM4[4063]<=26'd23466548;
ROM1[4064]<=26'd1976370; ROM2[4064]<=26'd11288227; ROM3[4064]<=26'd9748813; ROM4[4064]<=26'd23465029;
ROM1[4065]<=26'd1988226; ROM2[4065]<=26'd11289093; ROM3[4065]<=26'd9742954; ROM4[4065]<=26'd23464364;
ROM1[4066]<=26'd2001516; ROM2[4066]<=26'd11293480; ROM3[4066]<=26'd9740890; ROM4[4066]<=26'd23467829;
ROM1[4067]<=26'd1996007; ROM2[4067]<=26'd11292054; ROM3[4067]<=26'd9738762; ROM4[4067]<=26'd23466853;
ROM1[4068]<=26'd1985472; ROM2[4068]<=26'd11289033; ROM3[4068]<=26'd9738189; ROM4[4068]<=26'd23464408;
ROM1[4069]<=26'd1982099; ROM2[4069]<=26'd11290885; ROM3[4069]<=26'd9743546; ROM4[4069]<=26'd23465989;
ROM1[4070]<=26'd1978759; ROM2[4070]<=26'd11292488; ROM3[4070]<=26'd9750038; ROM4[4070]<=26'd23468490;
ROM1[4071]<=26'd1976038; ROM2[4071]<=26'd11291940; ROM3[4071]<=26'd9753258; ROM4[4071]<=26'd23469122;
ROM1[4072]<=26'd1981868; ROM2[4072]<=26'd11294797; ROM3[4072]<=26'd9755156; ROM4[4072]<=26'd23470755;
ROM1[4073]<=26'd1994073; ROM2[4073]<=26'd11296778; ROM3[4073]<=26'd9751693; ROM4[4073]<=26'd23471381;
ROM1[4074]<=26'd2004619; ROM2[4074]<=26'd11296034; ROM3[4074]<=26'd9745777; ROM4[4074]<=26'd23470925;
ROM1[4075]<=26'd2008107; ROM2[4075]<=26'd11299207; ROM3[4075]<=26'd9746527; ROM4[4075]<=26'd23474059;
ROM1[4076]<=26'd2000589; ROM2[4076]<=26'd11298320; ROM3[4076]<=26'd9747688; ROM4[4076]<=26'd23474890;
ROM1[4077]<=26'd1988490; ROM2[4077]<=26'd11293402; ROM3[4077]<=26'd9747622; ROM4[4077]<=26'd23473716;
ROM1[4078]<=26'd1980953; ROM2[4078]<=26'd11290771; ROM3[4078]<=26'd9746978; ROM4[4078]<=26'd23471636;
ROM1[4079]<=26'd1974967; ROM2[4079]<=26'd11289523; ROM3[4079]<=26'd9747808; ROM4[4079]<=26'd23470259;
ROM1[4080]<=26'd1982275; ROM2[4080]<=26'd11295507; ROM3[4080]<=26'd9752216; ROM4[4080]<=26'd23475248;
ROM1[4081]<=26'd1991444; ROM2[4081]<=26'd11298322; ROM3[4081]<=26'd9750146; ROM4[4081]<=26'd23475421;
ROM1[4082]<=26'd1997508; ROM2[4082]<=26'd11292083; ROM3[4082]<=26'd9737328; ROM4[4082]<=26'd23468419;
ROM1[4083]<=26'd1999877; ROM2[4083]<=26'd11289130; ROM3[4083]<=26'd9732221; ROM4[4083]<=26'd23465533;
ROM1[4084]<=26'd1993459; ROM2[4084]<=26'd11288774; ROM3[4084]<=26'd9736716; ROM4[4084]<=26'd23467667;
ROM1[4085]<=26'd1996204; ROM2[4085]<=26'd11297659; ROM3[4085]<=26'd9750061; ROM4[4085]<=26'd23477987;
ROM1[4086]<=26'd1994513; ROM2[4086]<=26'd11300901; ROM3[4086]<=26'd9756991; ROM4[4086]<=26'd23481698;
ROM1[4087]<=26'd1982135; ROM2[4087]<=26'd11293771; ROM3[4087]<=26'd9754884; ROM4[4087]<=26'd23476221;
ROM1[4088]<=26'd1979853; ROM2[4088]<=26'd11293376; ROM3[4088]<=26'd9754104; ROM4[4088]<=26'd23474346;
ROM1[4089]<=26'd1981742; ROM2[4089]<=26'd11290160; ROM3[4089]<=26'd9750480; ROM4[4089]<=26'd23470221;
ROM1[4090]<=26'd1992274; ROM2[4090]<=26'd11291376; ROM3[4090]<=26'd9748772; ROM4[4090]<=26'd23470552;
ROM1[4091]<=26'd2006398; ROM2[4091]<=26'd11298377; ROM3[4091]<=26'd9750448; ROM4[4091]<=26'd23476685;
ROM1[4092]<=26'd2005253; ROM2[4092]<=26'd11297332; ROM3[4092]<=26'd9752160; ROM4[4092]<=26'd23477605;
ROM1[4093]<=26'd1994286; ROM2[4093]<=26'd11292548; ROM3[4093]<=26'd9751120; ROM4[4093]<=26'd23473949;
ROM1[4094]<=26'd1992637; ROM2[4094]<=26'd11296751; ROM3[4094]<=26'd9760467; ROM4[4094]<=26'd23478677;
ROM1[4095]<=26'd1988060; ROM2[4095]<=26'd11297573; ROM3[4095]<=26'd9766379; ROM4[4095]<=26'd23481112;
ROM1[4096]<=26'd1974431; ROM2[4096]<=26'd11288621; ROM3[4096]<=26'd9761153; ROM4[4096]<=26'd23474334;
ROM1[4097]<=26'd1977208; ROM2[4097]<=26'd11287224; ROM3[4097]<=26'd9759765; ROM4[4097]<=26'd23474269;
ROM1[4098]<=26'd1991874; ROM2[4098]<=26'd11288228; ROM3[4098]<=26'd9756461; ROM4[4098]<=26'd23475374;
ROM1[4099]<=26'd2011204; ROM2[4099]<=26'd11296791; ROM3[4099]<=26'd9758953; ROM4[4099]<=26'd23482917;
ROM1[4100]<=26'd2009866; ROM2[4100]<=26'd11295079; ROM3[4100]<=26'd9757254; ROM4[4100]<=26'd23481631;
ROM1[4101]<=26'd1995848; ROM2[4101]<=26'd11287477; ROM3[4101]<=26'd9754817; ROM4[4101]<=26'd23474000;
ROM1[4102]<=26'd1990879; ROM2[4102]<=26'd11290526; ROM3[4102]<=26'd9760407; ROM4[4102]<=26'd23477196;
ROM1[4103]<=26'd1986527; ROM2[4103]<=26'd11290753; ROM3[4103]<=26'd9762129; ROM4[4103]<=26'd23477174;
ROM1[4104]<=26'd1984337; ROM2[4104]<=26'd11291675; ROM3[4104]<=26'd9765733; ROM4[4104]<=26'd23479484;
ROM1[4105]<=26'd1989014; ROM2[4105]<=26'd11294994; ROM3[4105]<=26'd9769757; ROM4[4105]<=26'd23484297;
ROM1[4106]<=26'd1996209; ROM2[4106]<=26'd11297131; ROM3[4106]<=26'd9768081; ROM4[4106]<=26'd23484228;
ROM1[4107]<=26'd2006361; ROM2[4107]<=26'd11298451; ROM3[4107]<=26'd9762099; ROM4[4107]<=26'd23483915;
ROM1[4108]<=26'd2016733; ROM2[4108]<=26'd11305393; ROM3[4108]<=26'd9766057; ROM4[4108]<=26'd23490100;
ROM1[4109]<=26'd2017204; ROM2[4109]<=26'd11310917; ROM3[4109]<=26'd9771230; ROM4[4109]<=26'd23495492;
ROM1[4110]<=26'd2006283; ROM2[4110]<=26'd11307059; ROM3[4110]<=26'd9768753; ROM4[4110]<=26'd23491157;
ROM1[4111]<=26'd1998853; ROM2[4111]<=26'd11303034; ROM3[4111]<=26'd9766284; ROM4[4111]<=26'd23486501;
ROM1[4112]<=26'd1991278; ROM2[4112]<=26'd11300517; ROM3[4112]<=26'd9766442; ROM4[4112]<=26'd23485193;
ROM1[4113]<=26'd1983033; ROM2[4113]<=26'd11294954; ROM3[4113]<=26'd9763360; ROM4[4113]<=26'd23479547;
ROM1[4114]<=26'd1987106; ROM2[4114]<=26'd11293776; ROM3[4114]<=26'd9760823; ROM4[4114]<=26'd23477394;
ROM1[4115]<=26'd2000256; ROM2[4115]<=26'd11295450; ROM3[4115]<=26'd9758238; ROM4[4115]<=26'd23479203;
ROM1[4116]<=26'd2007145; ROM2[4116]<=26'd11295393; ROM3[4116]<=26'd9754005; ROM4[4116]<=26'd23477570;
ROM1[4117]<=26'd2003163; ROM2[4117]<=26'd11295636; ROM3[4117]<=26'd9754108; ROM4[4117]<=26'd23477302;
ROM1[4118]<=26'd1995650; ROM2[4118]<=26'd11294384; ROM3[4118]<=26'd9754554; ROM4[4118]<=26'd23476960;
ROM1[4119]<=26'd1988098; ROM2[4119]<=26'd11290562; ROM3[4119]<=26'd9755992; ROM4[4119]<=26'd23475383;
ROM1[4120]<=26'd1980082; ROM2[4120]<=26'd11289204; ROM3[4120]<=26'd9756545; ROM4[4120]<=26'd23473580;
ROM1[4121]<=26'd1980495; ROM2[4121]<=26'd11292334; ROM3[4121]<=26'd9761217; ROM4[4121]<=26'd23478123;
ROM1[4122]<=26'd1986374; ROM2[4122]<=26'd11293898; ROM3[4122]<=26'd9762735; ROM4[4122]<=26'd23481749;
ROM1[4123]<=26'd1996107; ROM2[4123]<=26'd11293552; ROM3[4123]<=26'd9757436; ROM4[4123]<=26'd23479365;
ROM1[4124]<=26'd2008556; ROM2[4124]<=26'd11293563; ROM3[4124]<=26'd9753163; ROM4[4124]<=26'd23478563;
ROM1[4125]<=26'd2005086; ROM2[4125]<=26'd11290929; ROM3[4125]<=26'd9749944; ROM4[4125]<=26'd23476534;
ROM1[4126]<=26'd1996579; ROM2[4126]<=26'd11290876; ROM3[4126]<=26'd9751780; ROM4[4126]<=26'd23477101;
ROM1[4127]<=26'd1994456; ROM2[4127]<=26'd11294518; ROM3[4127]<=26'd9760038; ROM4[4127]<=26'd23481616;
ROM1[4128]<=26'd1990304; ROM2[4128]<=26'd11293918; ROM3[4128]<=26'd9762234; ROM4[4128]<=26'd23482019;
ROM1[4129]<=26'd1984573; ROM2[4129]<=26'd11293078; ROM3[4129]<=26'd9763661; ROM4[4129]<=26'd23481035;
ROM1[4130]<=26'd1985612; ROM2[4130]<=26'd11293800; ROM3[4130]<=26'd9764882; ROM4[4130]<=26'd23481661;
ROM1[4131]<=26'd1998270; ROM2[4131]<=26'd11299962; ROM3[4131]<=26'd9766213; ROM4[4131]<=26'd23487117;
ROM1[4132]<=26'd2012719; ROM2[4132]<=26'd11301868; ROM3[4132]<=26'd9761747; ROM4[4132]<=26'd23486032;
ROM1[4133]<=26'd2008034; ROM2[4133]<=26'd11292124; ROM3[4133]<=26'd9749701; ROM4[4133]<=26'd23474632;
ROM1[4134]<=26'd1998956; ROM2[4134]<=26'd11286522; ROM3[4134]<=26'd9750200; ROM4[4134]<=26'd23473299;
ROM1[4135]<=26'd1988333; ROM2[4135]<=26'd11283508; ROM3[4135]<=26'd9751355; ROM4[4135]<=26'd23470582;
ROM1[4136]<=26'd1983107; ROM2[4136]<=26'd11284476; ROM3[4136]<=26'd9755372; ROM4[4136]<=26'd23470849;
ROM1[4137]<=26'd1983325; ROM2[4137]<=26'd11290129; ROM3[4137]<=26'd9763897; ROM4[4137]<=26'd23477579;
ROM1[4138]<=26'd1979361; ROM2[4138]<=26'd11289539; ROM3[4138]<=26'd9761240; ROM4[4138]<=26'd23474495;
ROM1[4139]<=26'd1979354; ROM2[4139]<=26'd11285087; ROM3[4139]<=26'd9751194; ROM4[4139]<=26'd23466209;
ROM1[4140]<=26'd1988682; ROM2[4140]<=26'd11283583; ROM3[4140]<=26'd9742662; ROM4[4140]<=26'd23463431;
ROM1[4141]<=26'd1998922; ROM2[4141]<=26'd11286965; ROM3[4141]<=26'd9740435; ROM4[4141]<=26'd23466880;
ROM1[4142]<=26'd2006616; ROM2[4142]<=26'd11295384; ROM3[4142]<=26'd9747979; ROM4[4142]<=26'd23475106;
ROM1[4143]<=26'd2001539; ROM2[4143]<=26'd11297894; ROM3[4143]<=26'd9751694; ROM4[4143]<=26'd23477777;
ROM1[4144]<=26'd1990029; ROM2[4144]<=26'd11293944; ROM3[4144]<=26'd9751760; ROM4[4144]<=26'd23474722;
ROM1[4145]<=26'd1983090; ROM2[4145]<=26'd11291463; ROM3[4145]<=26'd9753920; ROM4[4145]<=26'd23473443;
ROM1[4146]<=26'd1975307; ROM2[4146]<=26'd11287137; ROM3[4146]<=26'd9752346; ROM4[4146]<=26'd23469914;
ROM1[4147]<=26'd1974174; ROM2[4147]<=26'd11283831; ROM3[4147]<=26'd9749537; ROM4[4147]<=26'd23467570;
ROM1[4148]<=26'd1984987; ROM2[4148]<=26'd11285900; ROM3[4148]<=26'd9744333; ROM4[4148]<=26'd23465787;
ROM1[4149]<=26'd1997171; ROM2[4149]<=26'd11288791; ROM3[4149]<=26'd9739015; ROM4[4149]<=26'd23465554;
ROM1[4150]<=26'd1996049; ROM2[4150]<=26'd11288324; ROM3[4150]<=26'd9738174; ROM4[4150]<=26'd23463499;
ROM1[4151]<=26'd1990735; ROM2[4151]<=26'd11286598; ROM3[4151]<=26'd9743701; ROM4[4151]<=26'd23464315;
ROM1[4152]<=26'd1985164; ROM2[4152]<=26'd11286304; ROM3[4152]<=26'd9749848; ROM4[4152]<=26'd23468017;
ROM1[4153]<=26'd1981187; ROM2[4153]<=26'd11286113; ROM3[4153]<=26'd9752827; ROM4[4153]<=26'd23468301;
ROM1[4154]<=26'd1976866; ROM2[4154]<=26'd11286716; ROM3[4154]<=26'd9753712; ROM4[4154]<=26'd23466968;
ROM1[4155]<=26'd1977499; ROM2[4155]<=26'd11288825; ROM3[4155]<=26'd9753827; ROM4[4155]<=26'd23468670;
ROM1[4156]<=26'd1988898; ROM2[4156]<=26'd11292086; ROM3[4156]<=26'd9754101; ROM4[4156]<=26'd23471562;
ROM1[4157]<=26'd2002024; ROM2[4157]<=26'd11294599; ROM3[4157]<=26'd9749499; ROM4[4157]<=26'd23471408;
ROM1[4158]<=26'd2002283; ROM2[4158]<=26'd11290365; ROM3[4158]<=26'd9745823; ROM4[4158]<=26'd23468319;
ROM1[4159]<=26'd1996564; ROM2[4159]<=26'd11288891; ROM3[4159]<=26'd9746707; ROM4[4159]<=26'd23466852;
ROM1[4160]<=26'd1992087; ROM2[4160]<=26'd11293012; ROM3[4160]<=26'd9752454; ROM4[4160]<=26'd23470845;
ROM1[4161]<=26'd1986272; ROM2[4161]<=26'd11292906; ROM3[4161]<=26'd9756129; ROM4[4161]<=26'd23471216;
ROM1[4162]<=26'd1974932; ROM2[4162]<=26'd11288048; ROM3[4162]<=26'd9754400; ROM4[4162]<=26'd23466157;
ROM1[4163]<=26'd1969093; ROM2[4163]<=26'd11283551; ROM3[4163]<=26'd9749565; ROM4[4163]<=26'd23461501;
ROM1[4164]<=26'd1972352; ROM2[4164]<=26'd11281283; ROM3[4164]<=26'd9744606; ROM4[4164]<=26'd23458383;
ROM1[4165]<=26'd1987658; ROM2[4165]<=26'd11286061; ROM3[4165]<=26'd9742395; ROM4[4165]<=26'd23460768;
ROM1[4166]<=26'd1999010; ROM2[4166]<=26'd11291097; ROM3[4166]<=26'd9740812; ROM4[4166]<=26'd23464805;
ROM1[4167]<=26'd1994283; ROM2[4167]<=26'd11290110; ROM3[4167]<=26'd9740966; ROM4[4167]<=26'd23463793;
ROM1[4168]<=26'd1983630; ROM2[4168]<=26'd11286499; ROM3[4168]<=26'd9740254; ROM4[4168]<=26'd23461458;
ROM1[4169]<=26'd1975282; ROM2[4169]<=26'd11282815; ROM3[4169]<=26'd9741238; ROM4[4169]<=26'd23460101;
ROM1[4170]<=26'd1972025; ROM2[4170]<=26'd11283098; ROM3[4170]<=26'd9745951; ROM4[4170]<=26'd23462090;
ROM1[4171]<=26'd1970130; ROM2[4171]<=26'd11283482; ROM3[4171]<=26'd9748047; ROM4[4171]<=26'd23462384;
ROM1[4172]<=26'd1973954; ROM2[4172]<=26'd11284600; ROM3[4172]<=26'd9747061; ROM4[4172]<=26'd23462714;
ROM1[4173]<=26'd1984979; ROM2[4173]<=26'd11286640; ROM3[4173]<=26'd9743321; ROM4[4173]<=26'd23462360;
ROM1[4174]<=26'd1996848; ROM2[4174]<=26'd11286243; ROM3[4174]<=26'd9739177; ROM4[4174]<=26'd23462217;
ROM1[4175]<=26'd1999439; ROM2[4175]<=26'd11287683; ROM3[4175]<=26'd9742039; ROM4[4175]<=26'd23467725;
ROM1[4176]<=26'd1992914; ROM2[4176]<=26'd11287569; ROM3[4176]<=26'd9746122; ROM4[4176]<=26'd23469539;
ROM1[4177]<=26'd1987817; ROM2[4177]<=26'd11287681; ROM3[4177]<=26'd9750492; ROM4[4177]<=26'd23470409;
ROM1[4178]<=26'd1985500; ROM2[4178]<=26'd11288860; ROM3[4178]<=26'd9753549; ROM4[4178]<=26'd23472502;
ROM1[4179]<=26'd1982574; ROM2[4179]<=26'd11291221; ROM3[4179]<=26'd9761550; ROM4[4179]<=26'd23476072;
ROM1[4180]<=26'd1990306; ROM2[4180]<=26'd11297785; ROM3[4180]<=26'd9770040; ROM4[4180]<=26'd23484053;
ROM1[4181]<=26'd1998870; ROM2[4181]<=26'd11298340; ROM3[4181]<=26'd9768244; ROM4[4181]<=26'd23485626;
ROM1[4182]<=26'd2003272; ROM2[4182]<=26'd11291093; ROM3[4182]<=26'd9756477; ROM4[4182]<=26'd23478925;
ROM1[4183]<=26'd2001571; ROM2[4183]<=26'd11286098; ROM3[4183]<=26'd9748833; ROM4[4183]<=26'd23473179;
ROM1[4184]<=26'd1992814; ROM2[4184]<=26'd11283753; ROM3[4184]<=26'd9750014; ROM4[4184]<=26'd23470918;
ROM1[4185]<=26'd1987671; ROM2[4185]<=26'd11285059; ROM3[4185]<=26'd9754286; ROM4[4185]<=26'd23472912;
ROM1[4186]<=26'd1991403; ROM2[4186]<=26'd11292885; ROM3[4186]<=26'd9765174; ROM4[4186]<=26'd23481910;
ROM1[4187]<=26'd1987145; ROM2[4187]<=26'd11294901; ROM3[4187]<=26'd9770650; ROM4[4187]<=26'd23484035;
ROM1[4188]<=26'd1983050; ROM2[4188]<=26'd11292091; ROM3[4188]<=26'd9769016; ROM4[4188]<=26'd23480936;
ROM1[4189]<=26'd1986920; ROM2[4189]<=26'd11288637; ROM3[4189]<=26'd9763804; ROM4[4189]<=26'd23478858;
ROM1[4190]<=26'd1997664; ROM2[4190]<=26'd11283860; ROM3[4190]<=26'd9755592; ROM4[4190]<=26'd23474740;
ROM1[4191]<=26'd2006609; ROM2[4191]<=26'd11277928; ROM3[4191]<=26'd9748917; ROM4[4191]<=26'd23472883;
ROM1[4192]<=26'd2000507; ROM2[4192]<=26'd11269459; ROM3[4192]<=26'd9744036; ROM4[4192]<=26'd23469784;
ROM1[4193]<=26'd1990295; ROM2[4193]<=26'd11264319; ROM3[4193]<=26'd9745790; ROM4[4193]<=26'd23468918;
ROM1[4194]<=26'd1983213; ROM2[4194]<=26'd11262542; ROM3[4194]<=26'd9750073; ROM4[4194]<=26'd23471059;
ROM1[4195]<=26'd1976366; ROM2[4195]<=26'd11260581; ROM3[4195]<=26'd9750096; ROM4[4195]<=26'd23469910;
ROM1[4196]<=26'd1975554; ROM2[4196]<=26'd11260733; ROM3[4196]<=26'd9750775; ROM4[4196]<=26'd23469909;
ROM1[4197]<=26'd1979382; ROM2[4197]<=26'd11260990; ROM3[4197]<=26'd9752093; ROM4[4197]<=26'd23471586;
ROM1[4198]<=26'd1986727; ROM2[4198]<=26'd11260667; ROM3[4198]<=26'd9747718; ROM4[4198]<=26'd23470177;
ROM1[4199]<=26'd1999461; ROM2[4199]<=26'd11262831; ROM3[4199]<=26'd9743380; ROM4[4199]<=26'd23471621;
ROM1[4200]<=26'd2002780; ROM2[4200]<=26'd11264750; ROM3[4200]<=26'd9746721; ROM4[4200]<=26'd23474134;
ROM1[4201]<=26'd1997644; ROM2[4201]<=26'd11263990; ROM3[4201]<=26'd9750033; ROM4[4201]<=26'd23475749;
ROM1[4202]<=26'd1991283; ROM2[4202]<=26'd11266621; ROM3[4202]<=26'd9755940; ROM4[4202]<=26'd23477726;
ROM1[4203]<=26'd1984462; ROM2[4203]<=26'd11266097; ROM3[4203]<=26'd9757087; ROM4[4203]<=26'd23476125;
ROM1[4204]<=26'd1977456; ROM2[4204]<=26'd11264003; ROM3[4204]<=26'd9756628; ROM4[4204]<=26'd23474137;
ROM1[4205]<=26'd1977595; ROM2[4205]<=26'd11263194; ROM3[4205]<=26'd9755834; ROM4[4205]<=26'd23471193;
ROM1[4206]<=26'd1986166; ROM2[4206]<=26'd11264037; ROM3[4206]<=26'd9751280; ROM4[4206]<=26'd23470154;
ROM1[4207]<=26'd2002462; ROM2[4207]<=26'd11270732; ROM3[4207]<=26'd9750776; ROM4[4207]<=26'd23476330;
ROM1[4208]<=26'd2005663; ROM2[4208]<=26'd11272662; ROM3[4208]<=26'd9749286; ROM4[4208]<=26'd23476802;
ROM1[4209]<=26'd1996704; ROM2[4209]<=26'd11269562; ROM3[4209]<=26'd9747133; ROM4[4209]<=26'd23473075;
ROM1[4210]<=26'd1990781; ROM2[4210]<=26'd11269473; ROM3[4210]<=26'd9749237; ROM4[4210]<=26'd23473272;
ROM1[4211]<=26'd1985981; ROM2[4211]<=26'd11268230; ROM3[4211]<=26'd9751436; ROM4[4211]<=26'd23470696;
ROM1[4212]<=26'd1979947; ROM2[4212]<=26'd11267684; ROM3[4212]<=26'd9753533; ROM4[4212]<=26'd23471456;
ROM1[4213]<=26'd1983217; ROM2[4213]<=26'd11275560; ROM3[4213]<=26'd9760034; ROM4[4213]<=26'd23479362;
ROM1[4214]<=26'd1991922; ROM2[4214]<=26'd11279264; ROM3[4214]<=26'd9761710; ROM4[4214]<=26'd23483136;
ROM1[4215]<=26'd2003767; ROM2[4215]<=26'd11279726; ROM3[4215]<=26'd9755716; ROM4[4215]<=26'd23482101;
ROM1[4216]<=26'd2013099; ROM2[4216]<=26'd11281075; ROM3[4216]<=26'd9751867; ROM4[4216]<=26'd23481186;
ROM1[4217]<=26'd2003521; ROM2[4217]<=26'd11275287; ROM3[4217]<=26'd9747486; ROM4[4217]<=26'd23476004;
ROM1[4218]<=26'd1989792; ROM2[4218]<=26'd11269653; ROM3[4218]<=26'd9743374; ROM4[4218]<=26'd23470449;
ROM1[4219]<=26'd1984434; ROM2[4219]<=26'd11268993; ROM3[4219]<=26'd9745655; ROM4[4219]<=26'd23470711;
ROM1[4220]<=26'd1977819; ROM2[4220]<=26'd11266467; ROM3[4220]<=26'd9749004; ROM4[4220]<=26'd23470864;
ROM1[4221]<=26'd1974482; ROM2[4221]<=26'd11264613; ROM3[4221]<=26'd9751553; ROM4[4221]<=26'd23471594;
ROM1[4222]<=26'd1979381; ROM2[4222]<=26'd11266443; ROM3[4222]<=26'd9752476; ROM4[4222]<=26'd23472710;
ROM1[4223]<=26'd1994837; ROM2[4223]<=26'd11273902; ROM3[4223]<=26'd9755814; ROM4[4223]<=26'd23479432;
ROM1[4224]<=26'd2005671; ROM2[4224]<=26'd11275565; ROM3[4224]<=26'd9751210; ROM4[4224]<=26'd23479180;
ROM1[4225]<=26'd1997804; ROM2[4225]<=26'd11266807; ROM3[4225]<=26'd9742393; ROM4[4225]<=26'd23471500;
ROM1[4226]<=26'd1988891; ROM2[4226]<=26'd11261566; ROM3[4226]<=26'd9745078; ROM4[4226]<=26'd23470363;
ROM1[4227]<=26'd1981914; ROM2[4227]<=26'd11259960; ROM3[4227]<=26'd9749359; ROM4[4227]<=26'd23471216;
ROM1[4228]<=26'd1980149; ROM2[4228]<=26'd11262958; ROM3[4228]<=26'd9753483; ROM4[4228]<=26'd23475611;
ROM1[4229]<=26'd1973012; ROM2[4229]<=26'd11261386; ROM3[4229]<=26'd9753968; ROM4[4229]<=26'd23473298;
ROM1[4230]<=26'd1977476; ROM2[4230]<=26'd11265332; ROM3[4230]<=26'd9759174; ROM4[4230]<=26'd23476563;
ROM1[4231]<=26'd1992488; ROM2[4231]<=26'd11273431; ROM3[4231]<=26'd9765932; ROM4[4231]<=26'd23483675;
ROM1[4232]<=26'd1998406; ROM2[4232]<=26'd11266469; ROM3[4232]<=26'd9754931; ROM4[4232]<=26'd23478093;
ROM1[4233]<=26'd2001508; ROM2[4233]<=26'd11264648; ROM3[4233]<=26'd9749745; ROM4[4233]<=26'd23475093;
ROM1[4234]<=26'd1993627; ROM2[4234]<=26'd11261900; ROM3[4234]<=26'd9746651; ROM4[4234]<=26'd23471616;
ROM1[4235]<=26'd1979974; ROM2[4235]<=26'd11253581; ROM3[4235]<=26'd9741706; ROM4[4235]<=26'd23464866;
ROM1[4236]<=26'd1976885; ROM2[4236]<=26'd11254619; ROM3[4236]<=26'd9745918; ROM4[4236]<=26'd23466412;
ROM1[4237]<=26'd1976111; ROM2[4237]<=26'd11258760; ROM3[4237]<=26'd9753906; ROM4[4237]<=26'd23470341;
ROM1[4238]<=26'd1979159; ROM2[4238]<=26'd11262141; ROM3[4238]<=26'd9757096; ROM4[4238]<=26'd23474161;
ROM1[4239]<=26'd1985810; ROM2[4239]<=26'd11263418; ROM3[4239]<=26'd9752248; ROM4[4239]<=26'd23473783;
ROM1[4240]<=26'd1997276; ROM2[4240]<=26'd11266073; ROM3[4240]<=26'd9748683; ROM4[4240]<=26'd23473227;
ROM1[4241]<=26'd2007924; ROM2[4241]<=26'd11271463; ROM3[4241]<=26'd9748892; ROM4[4241]<=26'd23478419;
ROM1[4242]<=26'd2004882; ROM2[4242]<=26'd11273361; ROM3[4242]<=26'd9750200; ROM4[4242]<=26'd23478952;
ROM1[4243]<=26'd1990011; ROM2[4243]<=26'd11266005; ROM3[4243]<=26'd9746782; ROM4[4243]<=26'd23471690;
ROM1[4244]<=26'd1979768; ROM2[4244]<=26'd11261071; ROM3[4244]<=26'd9745616; ROM4[4244]<=26'd23467295;
ROM1[4245]<=26'd1977237; ROM2[4245]<=26'd11262185; ROM3[4245]<=26'd9749044; ROM4[4245]<=26'd23469037;
ROM1[4246]<=26'd1972692; ROM2[4246]<=26'd11261863; ROM3[4246]<=26'd9748354; ROM4[4246]<=26'd23468805;
ROM1[4247]<=26'd1973967; ROM2[4247]<=26'd11262463; ROM3[4247]<=26'd9747744; ROM4[4247]<=26'd23469126;
ROM1[4248]<=26'd1986743; ROM2[4248]<=26'd11264075; ROM3[4248]<=26'd9745382; ROM4[4248]<=26'd23470136;
ROM1[4249]<=26'd2001787; ROM2[4249]<=26'd11269021; ROM3[4249]<=26'd9744417; ROM4[4249]<=26'd23473387;
ROM1[4250]<=26'd2003647; ROM2[4250]<=26'd11272199; ROM3[4250]<=26'd9746462; ROM4[4250]<=26'd23475465;
ROM1[4251]<=26'd1993718; ROM2[4251]<=26'd11267924; ROM3[4251]<=26'd9745132; ROM4[4251]<=26'd23471075;
ROM1[4252]<=26'd1987628; ROM2[4252]<=26'd11267515; ROM3[4252]<=26'd9749774; ROM4[4252]<=26'd23471331;
ROM1[4253]<=26'd1982841; ROM2[4253]<=26'd11267204; ROM3[4253]<=26'd9754144; ROM4[4253]<=26'd23471606;
ROM1[4254]<=26'd1977323; ROM2[4254]<=26'd11265931; ROM3[4254]<=26'd9758128; ROM4[4254]<=26'd23471334;
ROM1[4255]<=26'd1981230; ROM2[4255]<=26'd11269298; ROM3[4255]<=26'd9761797; ROM4[4255]<=26'd23475626;
ROM1[4256]<=26'd1990514; ROM2[4256]<=26'd11270513; ROM3[4256]<=26'd9756742; ROM4[4256]<=26'd23474455;
ROM1[4257]<=26'd2002235; ROM2[4257]<=26'd11269733; ROM3[4257]<=26'd9749335; ROM4[4257]<=26'd23472267;
ROM1[4258]<=26'd2006985; ROM2[4258]<=26'd11269707; ROM3[4258]<=26'd9748251; ROM4[4258]<=26'd23473483;
ROM1[4259]<=26'd2003099; ROM2[4259]<=26'd11270644; ROM3[4259]<=26'd9750897; ROM4[4259]<=26'd23474776;
ROM1[4260]<=26'd1991870; ROM2[4260]<=26'd11266000; ROM3[4260]<=26'd9751408; ROM4[4260]<=26'd23471854;
ROM1[4261]<=26'd1984723; ROM2[4261]<=26'd11262386; ROM3[4261]<=26'd9751033; ROM4[4261]<=26'd23470864;
ROM1[4262]<=26'd1975925; ROM2[4262]<=26'd11259886; ROM3[4262]<=26'd9750675; ROM4[4262]<=26'd23468976;
ROM1[4263]<=26'd1974543; ROM2[4263]<=26'd11260110; ROM3[4263]<=26'd9752708; ROM4[4263]<=26'd23469815;
ROM1[4264]<=26'd1990288; ROM2[4264]<=26'd11269442; ROM3[4264]<=26'd9759865; ROM4[4264]<=26'd23479017;
ROM1[4265]<=26'd2000556; ROM2[4265]<=26'd11267835; ROM3[4265]<=26'd9751641; ROM4[4265]<=26'd23475915;
ROM1[4266]<=26'd2001662; ROM2[4266]<=26'd11261287; ROM3[4266]<=26'd9740086; ROM4[4266]<=26'd23469654;
ROM1[4267]<=26'd1997380; ROM2[4267]<=26'd11259322; ROM3[4267]<=26'd9740473; ROM4[4267]<=26'd23469061;
ROM1[4268]<=26'd1987336; ROM2[4268]<=26'd11255135; ROM3[4268]<=26'd9742044; ROM4[4268]<=26'd23467134;
ROM1[4269]<=26'd1981729; ROM2[4269]<=26'd11254689; ROM3[4269]<=26'd9747012; ROM4[4269]<=26'd23467794;
ROM1[4270]<=26'd1977985; ROM2[4270]<=26'd11254287; ROM3[4270]<=26'd9751181; ROM4[4270]<=26'd23468111;
ROM1[4271]<=26'd1974208; ROM2[4271]<=26'd11253057; ROM3[4271]<=26'd9751626; ROM4[4271]<=26'd23468267;
ROM1[4272]<=26'd1976138; ROM2[4272]<=26'd11252050; ROM3[4272]<=26'd9749896; ROM4[4272]<=26'd23468560;
ROM1[4273]<=26'd1988493; ROM2[4273]<=26'd11253684; ROM3[4273]<=26'd9748872; ROM4[4273]<=26'd23470355;
ROM1[4274]<=26'd2002123; ROM2[4274]<=26'd11253482; ROM3[4274]<=26'd9746968; ROM4[4274]<=26'd23472549;
ROM1[4275]<=26'd2000423; ROM2[4275]<=26'd11249340; ROM3[4275]<=26'd9746896; ROM4[4275]<=26'd23472067;
ROM1[4276]<=26'd1992025; ROM2[4276]<=26'd11246411; ROM3[4276]<=26'd9749588; ROM4[4276]<=26'd23472282;
ROM1[4277]<=26'd1988102; ROM2[4277]<=26'd11248938; ROM3[4277]<=26'd9756348; ROM4[4277]<=26'd23476437;
ROM1[4278]<=26'd1985095; ROM2[4278]<=26'd11250770; ROM3[4278]<=26'd9759736; ROM4[4278]<=26'd23479752;
ROM1[4279]<=26'd1985204; ROM2[4279]<=26'd11254002; ROM3[4279]<=26'd9764236; ROM4[4279]<=26'd23482733;
ROM1[4280]<=26'd1988891; ROM2[4280]<=26'd11256803; ROM3[4280]<=26'd9765623; ROM4[4280]<=26'd23485289;
ROM1[4281]<=26'd1987866; ROM2[4281]<=26'd11245892; ROM3[4281]<=26'd9751806; ROM4[4281]<=26'd23474522;
ROM1[4282]<=26'd1996037; ROM2[4282]<=26'd11238938; ROM3[4282]<=26'd9741740; ROM4[4282]<=26'd23467758;
ROM1[4283]<=26'd1995173; ROM2[4283]<=26'd11234077; ROM3[4283]<=26'd9735177; ROM4[4283]<=26'd23463671;
ROM1[4284]<=26'd1984647; ROM2[4284]<=26'd11228735; ROM3[4284]<=26'd9730714; ROM4[4284]<=26'd23458116;
ROM1[4285]<=26'd1981495; ROM2[4285]<=26'd11229852; ROM3[4285]<=26'd9735130; ROM4[4285]<=26'd23460510;
ROM1[4286]<=26'd1980049; ROM2[4286]<=26'd11231421; ROM3[4286]<=26'd9739690; ROM4[4286]<=26'd23462466;
ROM1[4287]<=26'd1970721; ROM2[4287]<=26'd11227514; ROM3[4287]<=26'd9738394; ROM4[4287]<=26'd23460178;
ROM1[4288]<=26'd1965373; ROM2[4288]<=26'd11222979; ROM3[4288]<=26'd9735453; ROM4[4288]<=26'd23458289;
ROM1[4289]<=26'd1973505; ROM2[4289]<=26'd11225120; ROM3[4289]<=26'd9737981; ROM4[4289]<=26'd23462416;
ROM1[4290]<=26'd1989126; ROM2[4290]<=26'd11230865; ROM3[4290]<=26'd9737739; ROM4[4290]<=26'd23466650;
ROM1[4291]<=26'd2001542; ROM2[4291]<=26'd11235792; ROM3[4291]<=26'd9738677; ROM4[4291]<=26'd23471755;
ROM1[4292]<=26'd1998336; ROM2[4292]<=26'd11232785; ROM3[4292]<=26'd9740763; ROM4[4292]<=26'd23472407;
ROM1[4293]<=26'd1984565; ROM2[4293]<=26'd11225629; ROM3[4293]<=26'd9737628; ROM4[4293]<=26'd23467107;
ROM1[4294]<=26'd1974362; ROM2[4294]<=26'd11220661; ROM3[4294]<=26'd9737655; ROM4[4294]<=26'd23464146;
ROM1[4295]<=26'd1966235; ROM2[4295]<=26'd11216191; ROM3[4295]<=26'd9739400; ROM4[4295]<=26'd23461832;
ROM1[4296]<=26'd1966329; ROM2[4296]<=26'd11220043; ROM3[4296]<=26'd9744078; ROM4[4296]<=26'd23463978;
ROM1[4297]<=26'd1974476; ROM2[4297]<=26'd11226046; ROM3[4297]<=26'd9747565; ROM4[4297]<=26'd23467767;
ROM1[4298]<=26'd1985331; ROM2[4298]<=26'd11227823; ROM3[4298]<=26'd9744121; ROM4[4298]<=26'd23468947;
ROM1[4299]<=26'd2001409; ROM2[4299]<=26'd11232889; ROM3[4299]<=26'd9743109; ROM4[4299]<=26'd23473538;
ROM1[4300]<=26'd2001992; ROM2[4300]<=26'd11233168; ROM3[4300]<=26'd9743778; ROM4[4300]<=26'd23475448;
ROM1[4301]<=26'd1990698; ROM2[4301]<=26'd11229151; ROM3[4301]<=26'd9742875; ROM4[4301]<=26'd23472806;
ROM1[4302]<=26'd1983230; ROM2[4302]<=26'd11226582; ROM3[4302]<=26'd9746031; ROM4[4302]<=26'd23470683;
ROM1[4303]<=26'd1976778; ROM2[4303]<=26'd11225506; ROM3[4303]<=26'd9747144; ROM4[4303]<=26'd23468578;
ROM1[4304]<=26'd1968928; ROM2[4304]<=26'd11224325; ROM3[4304]<=26'd9747746; ROM4[4304]<=26'd23465353;
ROM1[4305]<=26'd1973765; ROM2[4305]<=26'd11227309; ROM3[4305]<=26'd9751477; ROM4[4305]<=26'd23468326;
ROM1[4306]<=26'd1985266; ROM2[4306]<=26'd11230781; ROM3[4306]<=26'd9751006; ROM4[4306]<=26'd23471896;
ROM1[4307]<=26'd1996870; ROM2[4307]<=26'd11230646; ROM3[4307]<=26'd9743553; ROM4[4307]<=26'd23469027;
ROM1[4308]<=26'd2003289; ROM2[4308]<=26'd11232798; ROM3[4308]<=26'd9743245; ROM4[4308]<=26'd23470985;
ROM1[4309]<=26'd1996224; ROM2[4309]<=26'd11231914; ROM3[4309]<=26'd9746189; ROM4[4309]<=26'd23471648;
ROM1[4310]<=26'd1988440; ROM2[4310]<=26'd11233209; ROM3[4310]<=26'd9749539; ROM4[4310]<=26'd23471527;
ROM1[4311]<=26'd1982079; ROM2[4311]<=26'd11233475; ROM3[4311]<=26'd9751354; ROM4[4311]<=26'd23471198;
ROM1[4312]<=26'd1968192; ROM2[4312]<=26'd11226140; ROM3[4312]<=26'd9747127; ROM4[4312]<=26'd23464562;
ROM1[4313]<=26'd1966095; ROM2[4313]<=26'd11225384; ROM3[4313]<=26'd9746986; ROM4[4313]<=26'd23463953;
ROM1[4314]<=26'd1970448; ROM2[4314]<=26'd11224219; ROM3[4314]<=26'd9743512; ROM4[4314]<=26'd23463790;
ROM1[4315]<=26'd1978678; ROM2[4315]<=26'd11220560; ROM3[4315]<=26'd9735075; ROM4[4315]<=26'd23459576;
ROM1[4316]<=26'd1987511; ROM2[4316]<=26'd11219461; ROM3[4316]<=26'd9732003; ROM4[4316]<=26'd23458048;
ROM1[4317]<=26'd1985247; ROM2[4317]<=26'd11221401; ROM3[4317]<=26'd9733242; ROM4[4317]<=26'd23459328;
ROM1[4318]<=26'd1977409; ROM2[4318]<=26'd11222986; ROM3[4318]<=26'd9737307; ROM4[4318]<=26'd23460515;
ROM1[4319]<=26'd1972461; ROM2[4319]<=26'd11221582; ROM3[4319]<=26'd9741047; ROM4[4319]<=26'd23460434;
ROM1[4320]<=26'd1970357; ROM2[4320]<=26'd11224927; ROM3[4320]<=26'd9746062; ROM4[4320]<=26'd23463541;
ROM1[4321]<=26'd1967307; ROM2[4321]<=26'd11226335; ROM3[4321]<=26'd9749795; ROM4[4321]<=26'd23464334;
ROM1[4322]<=26'd1972688; ROM2[4322]<=26'd11228608; ROM3[4322]<=26'd9749114; ROM4[4322]<=26'd23464816;
ROM1[4323]<=26'd1987973; ROM2[4323]<=26'd11235921; ROM3[4323]<=26'd9747458; ROM4[4323]<=26'd23468864;
ROM1[4324]<=26'd2001108; ROM2[4324]<=26'd11241304; ROM3[4324]<=26'd9745147; ROM4[4324]<=26'd23471962;
ROM1[4325]<=26'd2002403; ROM2[4325]<=26'd11241741; ROM3[4325]<=26'd9744437; ROM4[4325]<=26'd23472381;
ROM1[4326]<=26'd1993980; ROM2[4326]<=26'd11237738; ROM3[4326]<=26'd9744521; ROM4[4326]<=26'd23470473;
ROM1[4327]<=26'd1984642; ROM2[4327]<=26'd11236687; ROM3[4327]<=26'd9748152; ROM4[4327]<=26'd23470024;
ROM1[4328]<=26'd1979216; ROM2[4328]<=26'd11237723; ROM3[4328]<=26'd9750640; ROM4[4328]<=26'd23470568;
ROM1[4329]<=26'd1973510; ROM2[4329]<=26'd11235976; ROM3[4329]<=26'd9750997; ROM4[4329]<=26'd23468699;
ROM1[4330]<=26'd1976242; ROM2[4330]<=26'd11237626; ROM3[4330]<=26'd9752386; ROM4[4330]<=26'd23470513;
ROM1[4331]<=26'd1993272; ROM2[4331]<=26'd11244950; ROM3[4331]<=26'd9758226; ROM4[4331]<=26'd23478474;
ROM1[4332]<=26'd2009215; ROM2[4332]<=26'd11247660; ROM3[4332]<=26'd9756256; ROM4[4332]<=26'd23479853;
ROM1[4333]<=26'd2003846; ROM2[4333]<=26'd11240657; ROM3[4333]<=26'd9747454; ROM4[4333]<=26'd23472692;
ROM1[4334]<=26'd1993625; ROM2[4334]<=26'd11235901; ROM3[4334]<=26'd9745906; ROM4[4334]<=26'd23469140;
ROM1[4335]<=26'd1979554; ROM2[4335]<=26'd11228351; ROM3[4335]<=26'd9740100; ROM4[4335]<=26'd23462422;
ROM1[4336]<=26'd1974828; ROM2[4336]<=26'd11228969; ROM3[4336]<=26'd9742166; ROM4[4336]<=26'd23462650;
ROM1[4337]<=26'd1974098; ROM2[4337]<=26'd11234553; ROM3[4337]<=26'd9751396; ROM4[4337]<=26'd23468707;
ROM1[4338]<=26'd1969144; ROM2[4338]<=26'd11232614; ROM3[4338]<=26'd9749064; ROM4[4338]<=26'd23465522;
ROM1[4339]<=26'd1972842; ROM2[4339]<=26'd11230937; ROM3[4339]<=26'd9744020; ROM4[4339]<=26'd23462212;
ROM1[4340]<=26'd1986351; ROM2[4340]<=26'd11232284; ROM3[4340]<=26'd9739489; ROM4[4340]<=26'd23463441;
ROM1[4341]<=26'd2001201; ROM2[4341]<=26'd11239662; ROM3[4341]<=26'd9741406; ROM4[4341]<=26'd23469456;
ROM1[4342]<=26'd2002532; ROM2[4342]<=26'd11242522; ROM3[4342]<=26'd9745103; ROM4[4342]<=26'd23472131;
ROM1[4343]<=26'd1993633; ROM2[4343]<=26'd11239503; ROM3[4343]<=26'd9744775; ROM4[4343]<=26'd23469784;
ROM1[4344]<=26'd1983835; ROM2[4344]<=26'd11234000; ROM3[4344]<=26'd9743793; ROM4[4344]<=26'd23465909;
ROM1[4345]<=26'd1976348; ROM2[4345]<=26'd11231573; ROM3[4345]<=26'd9742616; ROM4[4345]<=26'd23462998;
ROM1[4346]<=26'd1970629; ROM2[4346]<=26'd11231067; ROM3[4346]<=26'd9743705; ROM4[4346]<=26'd23460918;
ROM1[4347]<=26'd1971906; ROM2[4347]<=26'd11231396; ROM3[4347]<=26'd9743403; ROM4[4347]<=26'd23459634;
ROM1[4348]<=26'd1984485; ROM2[4348]<=26'd11236999; ROM3[4348]<=26'd9741545; ROM4[4348]<=26'd23459984;
ROM1[4349]<=26'd1995711; ROM2[4349]<=26'd11237161; ROM3[4349]<=26'd9735330; ROM4[4349]<=26'd23459333;
ROM1[4350]<=26'd1995129; ROM2[4350]<=26'd11234774; ROM3[4350]<=26'd9734288; ROM4[4350]<=26'd23459575;
ROM1[4351]<=26'd1989420; ROM2[4351]<=26'd11235068; ROM3[4351]<=26'd9740044; ROM4[4351]<=26'd23461066;
ROM1[4352]<=26'd1981898; ROM2[4352]<=26'd11234724; ROM3[4352]<=26'd9743471; ROM4[4352]<=26'd23462044;
ROM1[4353]<=26'd1974714; ROM2[4353]<=26'd11233956; ROM3[4353]<=26'd9745350; ROM4[4353]<=26'd23461198;
ROM1[4354]<=26'd1971193; ROM2[4354]<=26'd11236748; ROM3[4354]<=26'd9750032; ROM4[4354]<=26'd23463051;
ROM1[4355]<=26'd1973968; ROM2[4355]<=26'd11238411; ROM3[4355]<=26'd9751109; ROM4[4355]<=26'd23464334;
ROM1[4356]<=26'd1980884; ROM2[4356]<=26'd11237552; ROM3[4356]<=26'd9745511; ROM4[4356]<=26'd23462624;
ROM1[4357]<=26'd1992651; ROM2[4357]<=26'd11238386; ROM3[4357]<=26'd9739066; ROM4[4357]<=26'd23461086;
ROM1[4358]<=26'd1995521; ROM2[4358]<=26'd11236460; ROM3[4358]<=26'd9735773; ROM4[4358]<=26'd23458242;
ROM1[4359]<=26'd1990626; ROM2[4359]<=26'd11235179; ROM3[4359]<=26'd9737970; ROM4[4359]<=26'd23458645;
ROM1[4360]<=26'd1987054; ROM2[4360]<=26'd11236504; ROM3[4360]<=26'd9742993; ROM4[4360]<=26'd23461925;
ROM1[4361]<=26'd1990090; ROM2[4361]<=26'd11245383; ROM3[4361]<=26'd9753105; ROM4[4361]<=26'd23470609;
ROM1[4362]<=26'd1986184; ROM2[4362]<=26'd11248964; ROM3[4362]<=26'd9756324; ROM4[4362]<=26'd23472672;
ROM1[4363]<=26'd1977721; ROM2[4363]<=26'd11243585; ROM3[4363]<=26'd9750517; ROM4[4363]<=26'd23465304;
ROM1[4364]<=26'd1982044; ROM2[4364]<=26'd11243232; ROM3[4364]<=26'd9748387; ROM4[4364]<=26'd23465520;
ROM1[4365]<=26'd1993213; ROM2[4365]<=26'd11242164; ROM3[4365]<=26'd9742195; ROM4[4365]<=26'd23465254;
ROM1[4366]<=26'd1998108; ROM2[4366]<=26'd11240441; ROM3[4366]<=26'd9737444; ROM4[4366]<=26'd23463488;
ROM1[4367]<=26'd1998818; ROM2[4367]<=26'd11244584; ROM3[4367]<=26'd9742867; ROM4[4367]<=26'd23467299;
ROM1[4368]<=26'd1995587; ROM2[4368]<=26'd11249066; ROM3[4368]<=26'd9751295; ROM4[4368]<=26'd23471229;
ROM1[4369]<=26'd1988775; ROM2[4369]<=26'd11247299; ROM3[4369]<=26'd9754619; ROM4[4369]<=26'd23470488;
ROM1[4370]<=26'd1982872; ROM2[4370]<=26'd11246138; ROM3[4370]<=26'd9756401; ROM4[4370]<=26'd23470565;
ROM1[4371]<=26'd1980144; ROM2[4371]<=26'd11247518; ROM3[4371]<=26'd9760533; ROM4[4371]<=26'd23473815;
ROM1[4372]<=26'd1980805; ROM2[4372]<=26'd11246916; ROM3[4372]<=26'd9758066; ROM4[4372]<=26'd23471680;
ROM1[4373]<=26'd1991438; ROM2[4373]<=26'd11248127; ROM3[4373]<=26'd9751921; ROM4[4373]<=26'd23469325;
ROM1[4374]<=26'd2003892; ROM2[4374]<=26'd11251226; ROM3[4374]<=26'd9748074; ROM4[4374]<=26'd23469981;
ROM1[4375]<=26'd2000209; ROM2[4375]<=26'd11247886; ROM3[4375]<=26'd9744210; ROM4[4375]<=26'd23467706;
ROM1[4376]<=26'd1989235; ROM2[4376]<=26'd11242785; ROM3[4376]<=26'd9741620; ROM4[4376]<=26'd23463404;
ROM1[4377]<=26'd1982542; ROM2[4377]<=26'd11243340; ROM3[4377]<=26'd9744839; ROM4[4377]<=26'd23463760;
ROM1[4378]<=26'd1978521; ROM2[4378]<=26'd11243997; ROM3[4378]<=26'd9747671; ROM4[4378]<=26'd23466187;
ROM1[4379]<=26'd1975176; ROM2[4379]<=26'd11246685; ROM3[4379]<=26'd9750118; ROM4[4379]<=26'd23466288;
ROM1[4380]<=26'd1976611; ROM2[4380]<=26'd11248363; ROM3[4380]<=26'd9750186; ROM4[4380]<=26'd23467035;
ROM1[4381]<=26'd1985093; ROM2[4381]<=26'd11249626; ROM3[4381]<=26'd9747241; ROM4[4381]<=26'd23467708;
ROM1[4382]<=26'd1998112; ROM2[4382]<=26'd11250991; ROM3[4382]<=26'd9742179; ROM4[4382]<=26'd23468067;
ROM1[4383]<=26'd2007224; ROM2[4383]<=26'd11255224; ROM3[4383]<=26'd9741051; ROM4[4383]<=26'd23471936;
ROM1[4384]<=26'd2006789; ROM2[4384]<=26'd11258282; ROM3[4384]<=26'd9745180; ROM4[4384]<=26'd23474837;
ROM1[4385]<=26'd2000074; ROM2[4385]<=26'd11257337; ROM3[4385]<=26'd9749160; ROM4[4385]<=26'd23475109;
ROM1[4386]<=26'd1991284; ROM2[4386]<=26'd11254428; ROM3[4386]<=26'd9747011; ROM4[4386]<=26'd23471733;
ROM1[4387]<=26'd1975764; ROM2[4387]<=26'd11244926; ROM3[4387]<=26'd9740239; ROM4[4387]<=26'd23462168;
ROM1[4388]<=26'd1971029; ROM2[4388]<=26'd11241993; ROM3[4388]<=26'd9738380; ROM4[4388]<=26'd23460416;
ROM1[4389]<=26'd1978686; ROM2[4389]<=26'd11244986; ROM3[4389]<=26'd9738497; ROM4[4389]<=26'd23463382;
ROM1[4390]<=26'd1994992; ROM2[4390]<=26'd11248792; ROM3[4390]<=26'd9737261; ROM4[4390]<=26'd23464632;
ROM1[4391]<=26'd2003973; ROM2[4391]<=26'd11253613; ROM3[4391]<=26'd9736930; ROM4[4391]<=26'd23468297;
ROM1[4392]<=26'd1996792; ROM2[4392]<=26'd11250783; ROM3[4392]<=26'd9733960; ROM4[4392]<=26'd23465747;
ROM1[4393]<=26'd1985309; ROM2[4393]<=26'd11244409; ROM3[4393]<=26'd9731181; ROM4[4393]<=26'd23459760;
ROM1[4394]<=26'd1979287; ROM2[4394]<=26'd11245090; ROM3[4394]<=26'd9735066; ROM4[4394]<=26'd23460943;
ROM1[4395]<=26'd1975360; ROM2[4395]<=26'd11246348; ROM3[4395]<=26'd9738584; ROM4[4395]<=26'd23461510;
ROM1[4396]<=26'd1972146; ROM2[4396]<=26'd11248237; ROM3[4396]<=26'd9741119; ROM4[4396]<=26'd23461972;
ROM1[4397]<=26'd1977582; ROM2[4397]<=26'd11251250; ROM3[4397]<=26'd9742587; ROM4[4397]<=26'd23464342;
ROM1[4398]<=26'd1990173; ROM2[4398]<=26'd11251576; ROM3[4398]<=26'd9739339; ROM4[4398]<=26'd23465014;
ROM1[4399]<=26'd2003627; ROM2[4399]<=26'd11253790; ROM3[4399]<=26'd9738310; ROM4[4399]<=26'd23467627;
ROM1[4400]<=26'd2004822; ROM2[4400]<=26'd11255394; ROM3[4400]<=26'd9741027; ROM4[4400]<=26'd23469906;
ROM1[4401]<=26'd1996925; ROM2[4401]<=26'd11254516; ROM3[4401]<=26'd9745023; ROM4[4401]<=26'd23470854;
ROM1[4402]<=26'd1987207; ROM2[4402]<=26'd11252990; ROM3[4402]<=26'd9748682; ROM4[4402]<=26'd23469363;
ROM1[4403]<=26'd1985225; ROM2[4403]<=26'd11254733; ROM3[4403]<=26'd9753616; ROM4[4403]<=26'd23471736;
ROM1[4404]<=26'd1983695; ROM2[4404]<=26'd11256894; ROM3[4404]<=26'd9756155; ROM4[4404]<=26'd23472728;
ROM1[4405]<=26'd1977243; ROM2[4405]<=26'd11250149; ROM3[4405]<=26'd9748313; ROM4[4405]<=26'd23464458;
ROM1[4406]<=26'd1978148; ROM2[4406]<=26'd11243096; ROM3[4406]<=26'd9737215; ROM4[4406]<=26'd23457989;
ROM1[4407]<=26'd1990290; ROM2[4407]<=26'd11246714; ROM3[4407]<=26'd9729703; ROM4[4407]<=26'd23457504;
ROM1[4408]<=26'd1993050; ROM2[4408]<=26'd11247886; ROM3[4408]<=26'd9728451; ROM4[4408]<=26'd23457386;
ROM1[4409]<=26'd1987827; ROM2[4409]<=26'd11248941; ROM3[4409]<=26'd9730268; ROM4[4409]<=26'd23458299;
ROM1[4410]<=26'd1985257; ROM2[4410]<=26'd11253495; ROM3[4410]<=26'd9737195; ROM4[4410]<=26'd23462466;
ROM1[4411]<=26'd1979999; ROM2[4411]<=26'd11254402; ROM3[4411]<=26'd9742918; ROM4[4411]<=26'd23465573;
ROM1[4412]<=26'd1970324; ROM2[4412]<=26'd11250228; ROM3[4412]<=26'd9741840; ROM4[4412]<=26'd23463508;
ROM1[4413]<=26'd1969821; ROM2[4413]<=26'd11249742; ROM3[4413]<=26'd9742212; ROM4[4413]<=26'd23462593;
ROM1[4414]<=26'd1975562; ROM2[4414]<=26'd11249918; ROM3[4414]<=26'd9739896; ROM4[4414]<=26'd23461512;
ROM1[4415]<=26'd1989372; ROM2[4415]<=26'd11250577; ROM3[4415]<=26'd9737493; ROM4[4415]<=26'd23462783;
ROM1[4416]<=26'd2004726; ROM2[4416]<=26'd11256903; ROM3[4416]<=26'd9742171; ROM4[4416]<=26'd23468917;
ROM1[4417]<=26'd2005571; ROM2[4417]<=26'd11263197; ROM3[4417]<=26'd9748216; ROM4[4417]<=26'd23475425;
ROM1[4418]<=26'd1996485; ROM2[4418]<=26'd11261356; ROM3[4418]<=26'd9749851; ROM4[4418]<=26'd23474219;
ROM1[4419]<=26'd1989584; ROM2[4419]<=26'd11259382; ROM3[4419]<=26'd9751085; ROM4[4419]<=26'd23472237;
ROM1[4420]<=26'd1978923; ROM2[4420]<=26'd11254342; ROM3[4420]<=26'd9748432; ROM4[4420]<=26'd23467995;
ROM1[4421]<=26'd1970503; ROM2[4421]<=26'd11248453; ROM3[4421]<=26'd9746702; ROM4[4421]<=26'd23463137;
ROM1[4422]<=26'd1977062; ROM2[4422]<=26'd11252360; ROM3[4422]<=26'd9749521; ROM4[4422]<=26'd23467196;
ROM1[4423]<=26'd1985711; ROM2[4423]<=26'd11251385; ROM3[4423]<=26'd9743957; ROM4[4423]<=26'd23464187;
ROM1[4424]<=26'd1994962; ROM2[4424]<=26'd11249938; ROM3[4424]<=26'd9738080; ROM4[4424]<=26'd23462534;
ROM1[4425]<=26'd1995654; ROM2[4425]<=26'd11250733; ROM3[4425]<=26'd9737233; ROM4[4425]<=26'd23463928;
ROM1[4426]<=26'd1988230; ROM2[4426]<=26'd11249465; ROM3[4426]<=26'd9738437; ROM4[4426]<=26'd23462858;
ROM1[4427]<=26'd1978575; ROM2[4427]<=26'd11248064; ROM3[4427]<=26'd9739891; ROM4[4427]<=26'd23462334;
ROM1[4428]<=26'd1972894; ROM2[4428]<=26'd11246802; ROM3[4428]<=26'd9742073; ROM4[4428]<=26'd23461042;
ROM1[4429]<=26'd1968028; ROM2[4429]<=26'd11246417; ROM3[4429]<=26'd9743225; ROM4[4429]<=26'd23459091;
ROM1[4430]<=26'd1966141; ROM2[4430]<=26'd11245462; ROM3[4430]<=26'd9740396; ROM4[4430]<=26'd23456515;
ROM1[4431]<=26'd1977049; ROM2[4431]<=26'd11246834; ROM3[4431]<=26'd9736386; ROM4[4431]<=26'd23456427;
ROM1[4432]<=26'd1993791; ROM2[4432]<=26'd11251268; ROM3[4432]<=26'd9733205; ROM4[4432]<=26'd23458660;
ROM1[4433]<=26'd1995939; ROM2[4433]<=26'd11251147; ROM3[4433]<=26'd9731583; ROM4[4433]<=26'd23458021;
ROM1[4434]<=26'd1992516; ROM2[4434]<=26'd11252411; ROM3[4434]<=26'd9734254; ROM4[4434]<=26'd23458208;
ROM1[4435]<=26'd1989134; ROM2[4435]<=26'd11255629; ROM3[4435]<=26'd9739993; ROM4[4435]<=26'd23459820;
ROM1[4436]<=26'd1981146; ROM2[4436]<=26'd11254193; ROM3[4436]<=26'd9739346; ROM4[4436]<=26'd23458104;
ROM1[4437]<=26'd1975135; ROM2[4437]<=26'd11252713; ROM3[4437]<=26'd9742121; ROM4[4437]<=26'd23459697;
ROM1[4438]<=26'd1983097; ROM2[4438]<=26'd11261224; ROM3[4438]<=26'd9751337; ROM4[4438]<=26'd23469448;
ROM1[4439]<=26'd1983226; ROM2[4439]<=26'd11257315; ROM3[4439]<=26'd9744578; ROM4[4439]<=26'd23464973;
ROM1[4440]<=26'd1982314; ROM2[4440]<=26'd11244142; ROM3[4440]<=26'd9727736; ROM4[4440]<=26'd23452194;
ROM1[4441]<=26'd1992265; ROM2[4441]<=26'd11247224; ROM3[4441]<=26'd9725864; ROM4[4441]<=26'd23455357;
ROM1[4442]<=26'd1989978; ROM2[4442]<=26'd11248710; ROM3[4442]<=26'd9729219; ROM4[4442]<=26'd23457200;
ROM1[4443]<=26'd1987866; ROM2[4443]<=26'd11252521; ROM3[4443]<=26'd9735148; ROM4[4443]<=26'd23460576;
ROM1[4444]<=26'd1988768; ROM2[4444]<=26'd11258081; ROM3[4444]<=26'd9743309; ROM4[4444]<=26'd23467000;
ROM1[4445]<=26'd1977385; ROM2[4445]<=26'd11250568; ROM3[4445]<=26'd9739936; ROM4[4445]<=26'd23460893;
ROM1[4446]<=26'd1969418; ROM2[4446]<=26'd11246484; ROM3[4446]<=26'd9737299; ROM4[4446]<=26'd23456430;
ROM1[4447]<=26'd1970720; ROM2[4447]<=26'd11246104; ROM3[4447]<=26'd9734715; ROM4[4447]<=26'd23455371;
ROM1[4448]<=26'd1982953; ROM2[4448]<=26'd11248805; ROM3[4448]<=26'd9732445; ROM4[4448]<=26'd23456382;
ROM1[4449]<=26'd1998412; ROM2[4449]<=26'd11254921; ROM3[4449]<=26'd9732296; ROM4[4449]<=26'd23459720;
ROM1[4450]<=26'd1999063; ROM2[4450]<=26'd11255719; ROM3[4450]<=26'd9733289; ROM4[4450]<=26'd23460554;
ROM1[4451]<=26'd1995552; ROM2[4451]<=26'd11258678; ROM3[4451]<=26'd9739506; ROM4[4451]<=26'd23464819;
ROM1[4452]<=26'd1989382; ROM2[4452]<=26'd11259973; ROM3[4452]<=26'd9743112; ROM4[4452]<=26'd23466029;
ROM1[4453]<=26'd1978003; ROM2[4453]<=26'd11251919; ROM3[4453]<=26'd9739279; ROM4[4453]<=26'd23460196;
ROM1[4454]<=26'd1967603; ROM2[4454]<=26'd11245748; ROM3[4454]<=26'd9735558; ROM4[4454]<=26'd23453973;
ROM1[4455]<=26'd1967134; ROM2[4455]<=26'd11244805; ROM3[4455]<=26'd9734090; ROM4[4455]<=26'd23451542;
ROM1[4456]<=26'd1973719; ROM2[4456]<=26'd11243776; ROM3[4456]<=26'd9729888; ROM4[4456]<=26'd23449624;
ROM1[4457]<=26'd1992173; ROM2[4457]<=26'd11250745; ROM3[4457]<=26'd9730130; ROM4[4457]<=26'd23454205;
ROM1[4458]<=26'd1997495; ROM2[4458]<=26'd11252549; ROM3[4458]<=26'd9729557; ROM4[4458]<=26'd23456035;
ROM1[4459]<=26'd1989686; ROM2[4459]<=26'd11249235; ROM3[4459]<=26'd9727512; ROM4[4459]<=26'd23454750;
ROM1[4460]<=26'd1985995; ROM2[4460]<=26'd11251461; ROM3[4460]<=26'd9732580; ROM4[4460]<=26'd23457629;
ROM1[4461]<=26'd1982144; ROM2[4461]<=26'd11252131; ROM3[4461]<=26'd9735638; ROM4[4461]<=26'd23456919;
ROM1[4462]<=26'd1981021; ROM2[4462]<=26'd11257319; ROM3[4462]<=26'd9742626; ROM4[4462]<=26'd23462509;
ROM1[4463]<=26'd1982842; ROM2[4463]<=26'd11258556; ROM3[4463]<=26'd9748330; ROM4[4463]<=26'd23466411;
ROM1[4464]<=26'd1988580; ROM2[4464]<=26'd11258328; ROM3[4464]<=26'd9747143; ROM4[4464]<=26'd23464881;
ROM1[4465]<=26'd1999829; ROM2[4465]<=26'd11259403; ROM3[4465]<=26'd9741370; ROM4[4465]<=26'd23464704;
ROM1[4466]<=26'd2003793; ROM2[4466]<=26'd11254414; ROM3[4466]<=26'd9734414; ROM4[4466]<=26'd23461144;
ROM1[4467]<=26'd1999984; ROM2[4467]<=26'd11252766; ROM3[4467]<=26'd9735159; ROM4[4467]<=26'd23460062;
ROM1[4468]<=26'd1991671; ROM2[4468]<=26'd11251927; ROM3[4468]<=26'd9738464; ROM4[4468]<=26'd23460179;
ROM1[4469]<=26'd1987035; ROM2[4469]<=26'd11251695; ROM3[4469]<=26'd9742423; ROM4[4469]<=26'd23461918;
ROM1[4470]<=26'd1979527; ROM2[4470]<=26'd11249572; ROM3[4470]<=26'd9743619; ROM4[4470]<=26'd23462133;
ROM1[4471]<=26'd1971290; ROM2[4471]<=26'd11245606; ROM3[4471]<=26'd9741841; ROM4[4471]<=26'd23458082;
ROM1[4472]<=26'd1977237; ROM2[4472]<=26'd11249568; ROM3[4472]<=26'd9742180; ROM4[4472]<=26'd23460073;
ROM1[4473]<=26'd1992328; ROM2[4473]<=26'd11256613; ROM3[4473]<=26'd9742719; ROM4[4473]<=26'd23465608;
ROM1[4474]<=26'd2001164; ROM2[4474]<=26'd11256149; ROM3[4474]<=26'd9737150; ROM4[4474]<=26'd23463480;
ROM1[4475]<=26'd1998295; ROM2[4475]<=26'd11252930; ROM3[4475]<=26'd9736873; ROM4[4475]<=26'd23461816;
ROM1[4476]<=26'd1993691; ROM2[4476]<=26'd11253114; ROM3[4476]<=26'd9743810; ROM4[4476]<=26'd23465079;
ROM1[4477]<=26'd1987667; ROM2[4477]<=26'd11252353; ROM3[4477]<=26'd9747493; ROM4[4477]<=26'd23465181;
ROM1[4478]<=26'd1980657; ROM2[4478]<=26'd11250491; ROM3[4478]<=26'd9749841; ROM4[4478]<=26'd23463978;
ROM1[4479]<=26'd1975519; ROM2[4479]<=26'd11248964; ROM3[4479]<=26'd9752679; ROM4[4479]<=26'd23463701;
ROM1[4480]<=26'd1978070; ROM2[4480]<=26'd11250174; ROM3[4480]<=26'd9753984; ROM4[4480]<=26'd23464668;
ROM1[4481]<=26'd1984408; ROM2[4481]<=26'd11249086; ROM3[4481]<=26'd9749786; ROM4[4481]<=26'd23463458;
ROM1[4482]<=26'd1996472; ROM2[4482]<=26'd11248647; ROM3[4482]<=26'd9744443; ROM4[4482]<=26'd23462296;
ROM1[4483]<=26'd2001434; ROM2[4483]<=26'd11248723; ROM3[4483]<=26'd9743399; ROM4[4483]<=26'd23462547;
ROM1[4484]<=26'd1996204; ROM2[4484]<=26'd11246342; ROM3[4484]<=26'd9744216; ROM4[4484]<=26'd23461947;
ROM1[4485]<=26'd1987260; ROM2[4485]<=26'd11243475; ROM3[4485]<=26'd9745815; ROM4[4485]<=26'd23459077;
ROM1[4486]<=26'd1982251; ROM2[4486]<=26'd11243731; ROM3[4486]<=26'd9747821; ROM4[4486]<=26'd23459343;
ROM1[4487]<=26'd1976891; ROM2[4487]<=26'd11247027; ROM3[4487]<=26'd9750911; ROM4[4487]<=26'd23462331;
ROM1[4488]<=26'd1973646; ROM2[4488]<=26'd11244746; ROM3[4488]<=26'd9749637; ROM4[4488]<=26'd23462000;
ROM1[4489]<=26'd1984548; ROM2[4489]<=26'd11249455; ROM3[4489]<=26'd9751823; ROM4[4489]<=26'd23466192;
ROM1[4490]<=26'd2002894; ROM2[4490]<=26'd11256581; ROM3[4490]<=26'd9753204; ROM4[4490]<=26'd23471064;
ROM1[4491]<=26'd2000670; ROM2[4491]<=26'd11245983; ROM3[4491]<=26'd9739427; ROM4[4491]<=26'd23460032;
ROM1[4492]<=26'd1991667; ROM2[4492]<=26'd11240949; ROM3[4492]<=26'd9734298; ROM4[4492]<=26'd23454396;
ROM1[4493]<=26'd1984279; ROM2[4493]<=26'd11239541; ROM3[4493]<=26'd9737585; ROM4[4493]<=26'd23455044;
ROM1[4494]<=26'd1976912; ROM2[4494]<=26'd11238622; ROM3[4494]<=26'd9741448; ROM4[4494]<=26'd23456150;
ROM1[4495]<=26'd1978774; ROM2[4495]<=26'd11248028; ROM3[4495]<=26'd9752265; ROM4[4495]<=26'd23465813;
ROM1[4496]<=26'd1981490; ROM2[4496]<=26'd11253802; ROM3[4496]<=26'd9758513; ROM4[4496]<=26'd23470921;
ROM1[4497]<=26'd1980323; ROM2[4497]<=26'd11248123; ROM3[4497]<=26'd9752211; ROM4[4497]<=26'd23466825;
ROM1[4498]<=26'd1989408; ROM2[4498]<=26'd11247079; ROM3[4498]<=26'd9743977; ROM4[4498]<=26'd23465190;
ROM1[4499]<=26'd2007539; ROM2[4499]<=26'd11255896; ROM3[4499]<=26'd9744507; ROM4[4499]<=26'd23471320;
ROM1[4500]<=26'd2005843; ROM2[4500]<=26'd11255493; ROM3[4500]<=26'd9743746; ROM4[4500]<=26'd23470951;
ROM1[4501]<=26'd1999650; ROM2[4501]<=26'd11256200; ROM3[4501]<=26'd9748618; ROM4[4501]<=26'd23473765;
ROM1[4502]<=26'd1995610; ROM2[4502]<=26'd11256781; ROM3[4502]<=26'd9757073; ROM4[4502]<=26'd23477730;
ROM1[4503]<=26'd1979618; ROM2[4503]<=26'd11244596; ROM3[4503]<=26'd9750680; ROM4[4503]<=26'd23469108;
ROM1[4504]<=26'd1970293; ROM2[4504]<=26'd11240135; ROM3[4504]<=26'd9749207; ROM4[4504]<=26'd23467226;
ROM1[4505]<=26'd1971956; ROM2[4505]<=26'd11242243; ROM3[4505]<=26'd9748801; ROM4[4505]<=26'd23466085;
ROM1[4506]<=26'd1978447; ROM2[4506]<=26'd11241250; ROM3[4506]<=26'd9740807; ROM4[4506]<=26'd23459755;
ROM1[4507]<=26'd1997669; ROM2[4507]<=26'd11248443; ROM3[4507]<=26'd9738980; ROM4[4507]<=26'd23462486;
ROM1[4508]<=26'd2004800; ROM2[4508]<=26'd11252791; ROM3[4508]<=26'd9742744; ROM4[4508]<=26'd23466643;
ROM1[4509]<=26'd2000278; ROM2[4509]<=26'd11252205; ROM3[4509]<=26'd9746006; ROM4[4509]<=26'd23468437;
ROM1[4510]<=26'd1991697; ROM2[4510]<=26'd11250476; ROM3[4510]<=26'd9747937; ROM4[4510]<=26'd23468173;
ROM1[4511]<=26'd1987277; ROM2[4511]<=26'd11250982; ROM3[4511]<=26'd9752654; ROM4[4511]<=26'd23469756;
ROM1[4512]<=26'd1981012; ROM2[4512]<=26'd11249479; ROM3[4512]<=26'd9753743; ROM4[4512]<=26'd23469123;
ROM1[4513]<=26'd1976417; ROM2[4513]<=26'd11245883; ROM3[4513]<=26'd9750748; ROM4[4513]<=26'd23464965;
ROM1[4514]<=26'd1981874; ROM2[4514]<=26'd11244454; ROM3[4514]<=26'd9746702; ROM4[4514]<=26'd23462811;
ROM1[4515]<=26'd1994630; ROM2[4515]<=26'd11245804; ROM3[4515]<=26'd9741029; ROM4[4515]<=26'd23463739;
ROM1[4516]<=26'd2002794; ROM2[4516]<=26'd11246619; ROM3[4516]<=26'd9738340; ROM4[4516]<=26'd23464223;
ROM1[4517]<=26'd1998628; ROM2[4517]<=26'd11246671; ROM3[4517]<=26'd9740311; ROM4[4517]<=26'd23464187;
ROM1[4518]<=26'd1993597; ROM2[4518]<=26'd11247273; ROM3[4518]<=26'd9744722; ROM4[4518]<=26'd23467021;
ROM1[4519]<=26'd1990790; ROM2[4519]<=26'd11246976; ROM3[4519]<=26'd9750680; ROM4[4519]<=26'd23470011;
ROM1[4520]<=26'd1988449; ROM2[4520]<=26'd11249367; ROM3[4520]<=26'd9755143; ROM4[4520]<=26'd23472003;
ROM1[4521]<=26'd1983749; ROM2[4521]<=26'd11247444; ROM3[4521]<=26'd9754410; ROM4[4521]<=26'd23471509;
ROM1[4522]<=26'd1984960; ROM2[4522]<=26'd11245278; ROM3[4522]<=26'd9750552; ROM4[4522]<=26'd23469155;
ROM1[4523]<=26'd1998246; ROM2[4523]<=26'd11249133; ROM3[4523]<=26'd9749291; ROM4[4523]<=26'd23470077;
ROM1[4524]<=26'd2011323; ROM2[4524]<=26'd11250914; ROM3[4524]<=26'd9748629; ROM4[4524]<=26'd23473150;
ROM1[4525]<=26'd2007834; ROM2[4525]<=26'd11247614; ROM3[4525]<=26'd9747544; ROM4[4525]<=26'd23471208;
ROM1[4526]<=26'd2001834; ROM2[4526]<=26'd11249384; ROM3[4526]<=26'd9752730; ROM4[4526]<=26'd23473819;
ROM1[4527]<=26'd1992644; ROM2[4527]<=26'd11245014; ROM3[4527]<=26'd9754640; ROM4[4527]<=26'd23472321;
ROM1[4528]<=26'd1979917; ROM2[4528]<=26'd11238929; ROM3[4528]<=26'd9751648; ROM4[4528]<=26'd23466453;
ROM1[4529]<=26'd1975699; ROM2[4529]<=26'd11241354; ROM3[4529]<=26'd9754798; ROM4[4529]<=26'd23468596;
ROM1[4530]<=26'd1976832; ROM2[4530]<=26'd11241125; ROM3[4530]<=26'd9754200; ROM4[4530]<=26'd23467621;
ROM1[4531]<=26'd1982680; ROM2[4531]<=26'd11239023; ROM3[4531]<=26'd9746085; ROM4[4531]<=26'd23463857;
ROM1[4532]<=26'd1995202; ROM2[4532]<=26'd11238983; ROM3[4532]<=26'd9739425; ROM4[4532]<=26'd23461913;
ROM1[4533]<=26'd1999942; ROM2[4533]<=26'd11240132; ROM3[4533]<=26'd9740056; ROM4[4533]<=26'd23463912;
ROM1[4534]<=26'd1993845; ROM2[4534]<=26'd11239911; ROM3[4534]<=26'd9741107; ROM4[4534]<=26'd23464770;
ROM1[4535]<=26'd1987598; ROM2[4535]<=26'd11242353; ROM3[4535]<=26'd9746816; ROM4[4535]<=26'd23468099;
ROM1[4536]<=26'd1989196; ROM2[4536]<=26'd11248086; ROM3[4536]<=26'd9756999; ROM4[4536]<=26'd23476616;
ROM1[4537]<=26'd1983218; ROM2[4537]<=26'd11247014; ROM3[4537]<=26'd9758848; ROM4[4537]<=26'd23475012;
ROM1[4538]<=26'd1978127; ROM2[4538]<=26'd11242618; ROM3[4538]<=26'd9754410; ROM4[4538]<=26'd23468614;
ROM1[4539]<=26'd1981153; ROM2[4539]<=26'd11237844; ROM3[4539]<=26'd9748845; ROM4[4539]<=26'd23464245;
ROM1[4540]<=26'd1984084; ROM2[4540]<=26'd11230954; ROM3[4540]<=26'd9735035; ROM4[4540]<=26'd23455195;
ROM1[4541]<=26'd1989429; ROM2[4541]<=26'd11229652; ROM3[4541]<=26'd9729158; ROM4[4541]<=26'd23452648;
ROM1[4542]<=26'd1988212; ROM2[4542]<=26'd11230621; ROM3[4542]<=26'd9736720; ROM4[4542]<=26'd23457475;
ROM1[4543]<=26'd1982199; ROM2[4543]<=26'd11231631; ROM3[4543]<=26'd9742098; ROM4[4543]<=26'd23459720;
ROM1[4544]<=26'd1976445; ROM2[4544]<=26'd11232222; ROM3[4544]<=26'd9745343; ROM4[4544]<=26'd23459163;
ROM1[4545]<=26'd1968680; ROM2[4545]<=26'd11230310; ROM3[4545]<=26'd9746195; ROM4[4545]<=26'd23458112;
ROM1[4546]<=26'd1965283; ROM2[4546]<=26'd11231505; ROM3[4546]<=26'd9747352; ROM4[4546]<=26'd23460404;
ROM1[4547]<=26'd1968090; ROM2[4547]<=26'd11231435; ROM3[4547]<=26'd9744255; ROM4[4547]<=26'd23458227;
ROM1[4548]<=26'd1978243; ROM2[4548]<=26'd11230559; ROM3[4548]<=26'd9737420; ROM4[4548]<=26'd23457042;
ROM1[4549]<=26'd1989764; ROM2[4549]<=26'd11232846; ROM3[4549]<=26'd9731693; ROM4[4549]<=26'd23458314;
ROM1[4550]<=26'd1987847; ROM2[4550]<=26'd11231231; ROM3[4550]<=26'd9727933; ROM4[4550]<=26'd23455752;
ROM1[4551]<=26'd1977554; ROM2[4551]<=26'd11227426; ROM3[4551]<=26'd9726001; ROM4[4551]<=26'd23451584;
ROM1[4552]<=26'd1976248; ROM2[4552]<=26'd11233420; ROM3[4552]<=26'd9732197; ROM4[4552]<=26'd23455786;
ROM1[4553]<=26'd1980615; ROM2[4553]<=26'd11242462; ROM3[4553]<=26'd9742479; ROM4[4553]<=26'd23462571;
ROM1[4554]<=26'd1970393; ROM2[4554]<=26'd11235766; ROM3[4554]<=26'd9739424; ROM4[4554]<=26'd23458638;
ROM1[4555]<=26'd1964721; ROM2[4555]<=26'd11228280; ROM3[4555]<=26'd9731900; ROM4[4555]<=26'd23452714;
ROM1[4556]<=26'd1972560; ROM2[4556]<=26'd11228792; ROM3[4556]<=26'd9728922; ROM4[4556]<=26'd23449531;
ROM1[4557]<=26'd1983204; ROM2[4557]<=26'd11229010; ROM3[4557]<=26'd9722650; ROM4[4557]<=26'd23447500;
ROM1[4558]<=26'd1988322; ROM2[4558]<=26'd11230337; ROM3[4558]<=26'd9723246; ROM4[4558]<=26'd23448565;
ROM1[4559]<=26'd1987789; ROM2[4559]<=26'd11233601; ROM3[4559]<=26'd9731186; ROM4[4559]<=26'd23454225;
ROM1[4560]<=26'd1978728; ROM2[4560]<=26'd11231065; ROM3[4560]<=26'd9733508; ROM4[4560]<=26'd23454478;
ROM1[4561]<=26'd1971763; ROM2[4561]<=26'd11227088; ROM3[4561]<=26'd9733833; ROM4[4561]<=26'd23453014;
ROM1[4562]<=26'd1970113; ROM2[4562]<=26'd11231207; ROM3[4562]<=26'd9739303; ROM4[4562]<=26'd23457094;
ROM1[4563]<=26'd1971372; ROM2[4563]<=26'd11233912; ROM3[4563]<=26'd9744115; ROM4[4563]<=26'd23460434;
ROM1[4564]<=26'd1974254; ROM2[4564]<=26'd11231076; ROM3[4564]<=26'd9739919; ROM4[4564]<=26'd23457518;
ROM1[4565]<=26'd1985175; ROM2[4565]<=26'd11230925; ROM3[4565]<=26'd9734557; ROM4[4565]<=26'd23456103;
ROM1[4566]<=26'd1996883; ROM2[4566]<=26'd11235407; ROM3[4566]<=26'd9736034; ROM4[4566]<=26'd23460246;
ROM1[4567]<=26'd1991628; ROM2[4567]<=26'd11234458; ROM3[4567]<=26'd9735795; ROM4[4567]<=26'd23458646;
ROM1[4568]<=26'd1981999; ROM2[4568]<=26'd11230183; ROM3[4568]<=26'd9735385; ROM4[4568]<=26'd23457299;
ROM1[4569]<=26'd1977241; ROM2[4569]<=26'd11230644; ROM3[4569]<=26'd9738720; ROM4[4569]<=26'd23459701;
ROM1[4570]<=26'd1968236; ROM2[4570]<=26'd11228447; ROM3[4570]<=26'd9739320; ROM4[4570]<=26'd23457219;
ROM1[4571]<=26'd1958879; ROM2[4571]<=26'd11221940; ROM3[4571]<=26'd9734583; ROM4[4571]<=26'd23450952;
ROM1[4572]<=26'd1962170; ROM2[4572]<=26'd11221876; ROM3[4572]<=26'd9735605; ROM4[4572]<=26'd23452784;
ROM1[4573]<=26'd1971413; ROM2[4573]<=26'd11220751; ROM3[4573]<=26'd9731858; ROM4[4573]<=26'd23453130;
ROM1[4574]<=26'd1979446; ROM2[4574]<=26'd11216234; ROM3[4574]<=26'd9722098; ROM4[4574]<=26'd23448074;
ROM1[4575]<=26'd1981826; ROM2[4575]<=26'd11218431; ROM3[4575]<=26'd9724393; ROM4[4575]<=26'd23450983;
ROM1[4576]<=26'd1974877; ROM2[4576]<=26'd11217206; ROM3[4576]<=26'd9727437; ROM4[4576]<=26'd23450418;
ROM1[4577]<=26'd1964267; ROM2[4577]<=26'd11212988; ROM3[4577]<=26'd9728103; ROM4[4577]<=26'd23445974;
ROM1[4578]<=26'd1960331; ROM2[4578]<=26'd11216339; ROM3[4578]<=26'd9734348; ROM4[4578]<=26'd23449142;
ROM1[4579]<=26'd1956658; ROM2[4579]<=26'd11218681; ROM3[4579]<=26'd9739482; ROM4[4579]<=26'd23452360;
ROM1[4580]<=26'd1954120; ROM2[4580]<=26'd11214931; ROM3[4580]<=26'd9733964; ROM4[4580]<=26'd23448307;
ROM1[4581]<=26'd1962081; ROM2[4581]<=26'd11213249; ROM3[4581]<=26'd9729730; ROM4[4581]<=26'd23445828;
ROM1[4582]<=26'd1973019; ROM2[4582]<=26'd11212801; ROM3[4582]<=26'd9722909; ROM4[4582]<=26'd23443045;
ROM1[4583]<=26'd1975673; ROM2[4583]<=26'd11213609; ROM3[4583]<=26'd9718559; ROM4[4583]<=26'd23441955;
ROM1[4584]<=26'd1973263; ROM2[4584]<=26'd11217243; ROM3[4584]<=26'd9722409; ROM4[4584]<=26'd23444713;
ROM1[4585]<=26'd1968700; ROM2[4585]<=26'd11219555; ROM3[4585]<=26'd9726894; ROM4[4585]<=26'd23446760;
ROM1[4586]<=26'd1964042; ROM2[4586]<=26'd11218383; ROM3[4586]<=26'd9728648; ROM4[4586]<=26'd23446273;
ROM1[4587]<=26'd1954220; ROM2[4587]<=26'd11212843; ROM3[4587]<=26'd9726380; ROM4[4587]<=26'd23442203;
ROM1[4588]<=26'd1952894; ROM2[4588]<=26'd11213360; ROM3[4588]<=26'd9726401; ROM4[4588]<=26'd23440141;
ROM1[4589]<=26'd1966063; ROM2[4589]<=26'd11220076; ROM3[4589]<=26'd9728567; ROM4[4589]<=26'd23445761;
ROM1[4590]<=26'd1977382; ROM2[4590]<=26'd11218453; ROM3[4590]<=26'd9721566; ROM4[4590]<=26'd23445541;
ROM1[4591]<=26'd1977424; ROM2[4591]<=26'd11212738; ROM3[4591]<=26'd9711403; ROM4[4591]<=26'd23439949;
ROM1[4592]<=26'd1973242; ROM2[4592]<=26'd11210940; ROM3[4592]<=26'd9713523; ROM4[4592]<=26'd23441098;
ROM1[4593]<=26'd1963884; ROM2[4593]<=26'd11206962; ROM3[4593]<=26'd9713451; ROM4[4593]<=26'd23438217;
ROM1[4594]<=26'd1959570; ROM2[4594]<=26'd11207696; ROM3[4594]<=26'd9717607; ROM4[4594]<=26'd23438390;
ROM1[4595]<=26'd1959398; ROM2[4595]<=26'd11213451; ROM3[4595]<=26'd9727112; ROM4[4595]<=26'd23443363;
ROM1[4596]<=26'd1959368; ROM2[4596]<=26'd11215140; ROM3[4596]<=26'd9731368; ROM4[4596]<=26'd23446781;
ROM1[4597]<=26'd1959990; ROM2[4597]<=26'd11212445; ROM3[4597]<=26'd9728827; ROM4[4597]<=26'd23445603;
ROM1[4598]<=26'd1970335; ROM2[4598]<=26'd11214890; ROM3[4598]<=26'd9724265; ROM4[4598]<=26'd23446258;
ROM1[4599]<=26'd1987169; ROM2[4599]<=26'd11221683; ROM3[4599]<=26'd9726108; ROM4[4599]<=26'd23452779;
ROM1[4600]<=26'd1987274; ROM2[4600]<=26'd11221454; ROM3[4600]<=26'd9726607; ROM4[4600]<=26'd23454659;
ROM1[4601]<=26'd1980379; ROM2[4601]<=26'd11221565; ROM3[4601]<=26'd9728261; ROM4[4601]<=26'd23454003;
ROM1[4602]<=26'd1971174; ROM2[4602]<=26'd11219690; ROM3[4602]<=26'd9729688; ROM4[4602]<=26'd23450784;
ROM1[4603]<=26'd1965542; ROM2[4603]<=26'd11216407; ROM3[4603]<=26'd9729235; ROM4[4603]<=26'd23449286;
ROM1[4604]<=26'd1956125; ROM2[4604]<=26'd11210789; ROM3[4604]<=26'd9725157; ROM4[4604]<=26'd23444745;
ROM1[4605]<=26'd1952318; ROM2[4605]<=26'd11207949; ROM3[4605]<=26'd9719796; ROM4[4605]<=26'd23440131;
ROM1[4606]<=26'd1960018; ROM2[4606]<=26'd11207881; ROM3[4606]<=26'd9716760; ROM4[4606]<=26'd23438739;
ROM1[4607]<=26'd1970872; ROM2[4607]<=26'd11206513; ROM3[4607]<=26'd9712094; ROM4[4607]<=26'd23436299;
ROM1[4608]<=26'd1975178; ROM2[4608]<=26'd11208131; ROM3[4608]<=26'd9713515; ROM4[4608]<=26'd23438904;
ROM1[4609]<=26'd1974601; ROM2[4609]<=26'd11211688; ROM3[4609]<=26'd9720745; ROM4[4609]<=26'd23444945;
ROM1[4610]<=26'd1966932; ROM2[4610]<=26'd11211652; ROM3[4610]<=26'd9723571; ROM4[4610]<=26'd23445392;
ROM1[4611]<=26'd1951092; ROM2[4611]<=26'd11203636; ROM3[4611]<=26'd9717545; ROM4[4611]<=26'd23435375;
ROM1[4612]<=26'd1940530; ROM2[4612]<=26'd11199450; ROM3[4612]<=26'd9713933; ROM4[4612]<=26'd23428796;
ROM1[4613]<=26'd1941697; ROM2[4613]<=26'd11200948; ROM3[4613]<=26'd9717803; ROM4[4613]<=26'd23431157;
ROM1[4614]<=26'd1952387; ROM2[4614]<=26'd11205904; ROM3[4614]<=26'd9722311; ROM4[4614]<=26'd23437224;
ROM1[4615]<=26'd1968186; ROM2[4615]<=26'd11209838; ROM3[4615]<=26'd9719742; ROM4[4615]<=26'd23440006;
ROM1[4616]<=26'd1974640; ROM2[4616]<=26'd11210463; ROM3[4616]<=26'd9716945; ROM4[4616]<=26'd23439296;
ROM1[4617]<=26'd1968499; ROM2[4617]<=26'd11207909; ROM3[4617]<=26'd9714101; ROM4[4617]<=26'd23436997;
ROM1[4618]<=26'd1961473; ROM2[4618]<=26'd11206023; ROM3[4618]<=26'd9714418; ROM4[4618]<=26'd23436819;
ROM1[4619]<=26'd1963292; ROM2[4619]<=26'd11213106; ROM3[4619]<=26'd9725805; ROM4[4619]<=26'd23445474;
ROM1[4620]<=26'd1968370; ROM2[4620]<=26'd11222760; ROM3[4620]<=26'd9738097; ROM4[4620]<=26'd23455094;
ROM1[4621]<=26'd1955933; ROM2[4621]<=26'd11213244; ROM3[4621]<=26'd9732357; ROM4[4621]<=26'd23446882;
ROM1[4622]<=26'd1951551; ROM2[4622]<=26'd11205237; ROM3[4622]<=26'd9721529; ROM4[4622]<=26'd23439226;
ROM1[4623]<=26'd1967394; ROM2[4623]<=26'd11210433; ROM3[4623]<=26'd9718912; ROM4[4623]<=26'd23443758;
ROM1[4624]<=26'd1980788; ROM2[4624]<=26'd11214704; ROM3[4624]<=26'd9717634; ROM4[4624]<=26'd23448075;
ROM1[4625]<=26'd1986080; ROM2[4625]<=26'd11220278; ROM3[4625]<=26'd9723894; ROM4[4625]<=26'd23455267;
ROM1[4626]<=26'd1982370; ROM2[4626]<=26'd11221945; ROM3[4626]<=26'd9730987; ROM4[4626]<=26'd23458423;
ROM1[4627]<=26'd1973938; ROM2[4627]<=26'd11220120; ROM3[4627]<=26'd9734839; ROM4[4627]<=26'd23458093;
ROM1[4628]<=26'd1966976; ROM2[4628]<=26'd11215936; ROM3[4628]<=26'd9734673; ROM4[4628]<=26'd23457490;
ROM1[4629]<=26'd1964004; ROM2[4629]<=26'd11217696; ROM3[4629]<=26'd9740165; ROM4[4629]<=26'd23458528;
ROM1[4630]<=26'd1970218; ROM2[4630]<=26'd11223876; ROM3[4630]<=26'd9747321; ROM4[4630]<=26'd23463336;
ROM1[4631]<=26'd1975921; ROM2[4631]<=26'd11221579; ROM3[4631]<=26'd9741023; ROM4[4631]<=26'd23459978;
ROM1[4632]<=26'd1983122; ROM2[4632]<=26'd11217006; ROM3[4632]<=26'd9732617; ROM4[4632]<=26'd23452878;
ROM1[4633]<=26'd1987251; ROM2[4633]<=26'd11218762; ROM3[4633]<=26'd9731536; ROM4[4633]<=26'd23453043;
ROM1[4634]<=26'd1987077; ROM2[4634]<=26'd11224530; ROM3[4634]<=26'd9739385; ROM4[4634]<=26'd23459766;
ROM1[4635]<=26'd1986136; ROM2[4635]<=26'd11230615; ROM3[4635]<=26'd9749588; ROM4[4635]<=26'd23467896;
ROM1[4636]<=26'd1974463; ROM2[4636]<=26'd11224845; ROM3[4636]<=26'd9744623; ROM4[4636]<=26'd23462227;
ROM1[4637]<=26'd1956964; ROM2[4637]<=26'd11213657; ROM3[4637]<=26'd9735836; ROM4[4637]<=26'd23451358;
ROM1[4638]<=26'd1952124; ROM2[4638]<=26'd11210786; ROM3[4638]<=26'd9731888; ROM4[4638]<=26'd23448252;
ROM1[4639]<=26'd1959342; ROM2[4639]<=26'd11210810; ROM3[4639]<=26'd9728768; ROM4[4639]<=26'd23448150;
ROM1[4640]<=26'd1978588; ROM2[4640]<=26'd11218832; ROM3[4640]<=26'd9730012; ROM4[4640]<=26'd23454507;
ROM1[4641]<=26'd1990140; ROM2[4641]<=26'd11222734; ROM3[4641]<=26'd9730451; ROM4[4641]<=26'd23459152;
ROM1[4642]<=26'd1982200; ROM2[4642]<=26'd11215652; ROM3[4642]<=26'd9727528; ROM4[4642]<=26'd23455499;
ROM1[4643]<=26'd1972122; ROM2[4643]<=26'd11212916; ROM3[4643]<=26'd9729781; ROM4[4643]<=26'd23452655;
ROM1[4644]<=26'd1968250; ROM2[4644]<=26'd11216548; ROM3[4644]<=26'd9735161; ROM4[4644]<=26'd23454527;
ROM1[4645]<=26'd1964140; ROM2[4645]<=26'd11218373; ROM3[4645]<=26'd9739110; ROM4[4645]<=26'd23456485;
ROM1[4646]<=26'd1958054; ROM2[4646]<=26'd11215884; ROM3[4646]<=26'd9739997; ROM4[4646]<=26'd23454309;
ROM1[4647]<=26'd1960896; ROM2[4647]<=26'd11216345; ROM3[4647]<=26'd9738868; ROM4[4647]<=26'd23454787;
ROM1[4648]<=26'd1975360; ROM2[4648]<=26'd11221029; ROM3[4648]<=26'd9739479; ROM4[4648]<=26'd23458299;
ROM1[4649]<=26'd1985842; ROM2[4649]<=26'd11221597; ROM3[4649]<=26'd9735103; ROM4[4649]<=26'd23459429;
ROM1[4650]<=26'd1982844; ROM2[4650]<=26'd11219998; ROM3[4650]<=26'd9731134; ROM4[4650]<=26'd23456976;
ROM1[4651]<=26'd1976100; ROM2[4651]<=26'd11218593; ROM3[4651]<=26'd9732781; ROM4[4651]<=26'd23455739;
ROM1[4652]<=26'd1966775; ROM2[4652]<=26'd11214561; ROM3[4652]<=26'd9734196; ROM4[4652]<=26'd23453296;
ROM1[4653]<=26'd1959313; ROM2[4653]<=26'd11211110; ROM3[4653]<=26'd9733418; ROM4[4653]<=26'd23450016;
ROM1[4654]<=26'd1955885; ROM2[4654]<=26'd11211280; ROM3[4654]<=26'd9734416; ROM4[4654]<=26'd23451559;
ROM1[4655]<=26'd1956014; ROM2[4655]<=26'd11211746; ROM3[4655]<=26'd9731554; ROM4[4655]<=26'd23450413;
ROM1[4656]<=26'd1963684; ROM2[4656]<=26'd11210582; ROM3[4656]<=26'd9724487; ROM4[4656]<=26'd23446086;
ROM1[4657]<=26'd1979910; ROM2[4657]<=26'd11212654; ROM3[4657]<=26'd9718358; ROM4[4657]<=26'd23446181;
ROM1[4658]<=26'd1985116; ROM2[4658]<=26'd11212031; ROM3[4658]<=26'd9716675; ROM4[4658]<=26'd23446535;
ROM1[4659]<=26'd1981137; ROM2[4659]<=26'd11212771; ROM3[4659]<=26'd9721401; ROM4[4659]<=26'd23447187;
ROM1[4660]<=26'd1972622; ROM2[4660]<=26'd11212336; ROM3[4660]<=26'd9725418; ROM4[4660]<=26'd23447837;
ROM1[4661]<=26'd1967262; ROM2[4661]<=26'd11210569; ROM3[4661]<=26'd9727932; ROM4[4661]<=26'd23447726;
ROM1[4662]<=26'd1963058; ROM2[4662]<=26'd11211180; ROM3[4662]<=26'd9731365; ROM4[4662]<=26'd23448835;
ROM1[4663]<=26'd1960070; ROM2[4663]<=26'd11210020; ROM3[4663]<=26'd9732499; ROM4[4663]<=26'd23448418;
ROM1[4664]<=26'd1965286; ROM2[4664]<=26'd11210145; ROM3[4664]<=26'd9727474; ROM4[4664]<=26'd23447053;
ROM1[4665]<=26'd1976196; ROM2[4665]<=26'd11211069; ROM3[4665]<=26'd9721171; ROM4[4665]<=26'd23445044;
ROM1[4666]<=26'd1984962; ROM2[4666]<=26'd11214456; ROM3[4666]<=26'd9721797; ROM4[4666]<=26'd23448266;
ROM1[4667]<=26'd1990682; ROM2[4667]<=26'd11222349; ROM3[4667]<=26'd9729272; ROM4[4667]<=26'd23457608;
ROM1[4668]<=26'd1988042; ROM2[4668]<=26'd11224151; ROM3[4668]<=26'd9736293; ROM4[4668]<=26'd23461659;
ROM1[4669]<=26'd1976185; ROM2[4669]<=26'd11218335; ROM3[4669]<=26'd9736324; ROM4[4669]<=26'd23458418;
ROM1[4670]<=26'd1970349; ROM2[4670]<=26'd11218134; ROM3[4670]<=26'd9737105; ROM4[4670]<=26'd23458030;
ROM1[4671]<=26'd1962009; ROM2[4671]<=26'd11211387; ROM3[4671]<=26'd9731452; ROM4[4671]<=26'd23452190;
ROM1[4672]<=26'd1958813; ROM2[4672]<=26'd11202966; ROM3[4672]<=26'd9722774; ROM4[4672]<=26'd23446259;
ROM1[4673]<=26'd1976103; ROM2[4673]<=26'd11211055; ROM3[4673]<=26'd9723199; ROM4[4673]<=26'd23452741;
ROM1[4674]<=26'd1986078; ROM2[4674]<=26'd11211388; ROM3[4674]<=26'd9718997; ROM4[4674]<=26'd23453243;
ROM1[4675]<=26'd1986598; ROM2[4675]<=26'd11211719; ROM3[4675]<=26'd9720881; ROM4[4675]<=26'd23454880;
ROM1[4676]<=26'd1988865; ROM2[4676]<=26'd11218958; ROM3[4676]<=26'd9731809; ROM4[4676]<=26'd23462334;
ROM1[4677]<=26'd1982066; ROM2[4677]<=26'd11218227; ROM3[4677]<=26'd9737652; ROM4[4677]<=26'd23463587;
ROM1[4678]<=26'd1974158; ROM2[4678]<=26'd11216115; ROM3[4678]<=26'd9739429; ROM4[4678]<=26'd23461800;
ROM1[4679]<=26'd1965887; ROM2[4679]<=26'd11212197; ROM3[4679]<=26'd9738095; ROM4[4679]<=26'd23458864;
ROM1[4680]<=26'd1964188; ROM2[4680]<=26'd11211464; ROM3[4680]<=26'd9737411; ROM4[4680]<=26'd23457365;
ROM1[4681]<=26'd1976532; ROM2[4681]<=26'd11215977; ROM3[4681]<=26'd9737567; ROM4[4681]<=26'd23459301;
ROM1[4682]<=26'd1993268; ROM2[4682]<=26'd11220298; ROM3[4682]<=26'd9735856; ROM4[4682]<=26'd23462633;
ROM1[4683]<=26'd1997877; ROM2[4683]<=26'd11221495; ROM3[4683]<=26'd9736175; ROM4[4683]<=26'd23463008;
ROM1[4684]<=26'd1989280; ROM2[4684]<=26'd11217628; ROM3[4684]<=26'd9734460; ROM4[4684]<=26'd23460523;
ROM1[4685]<=26'd1979756; ROM2[4685]<=26'd11215081; ROM3[4685]<=26'd9735984; ROM4[4685]<=26'd23460794;
ROM1[4686]<=26'd1976271; ROM2[4686]<=26'd11215272; ROM3[4686]<=26'd9741006; ROM4[4686]<=26'd23461772;
ROM1[4687]<=26'd1971817; ROM2[4687]<=26'd11215908; ROM3[4687]<=26'd9746058; ROM4[4687]<=26'd23464696;
ROM1[4688]<=26'd1975616; ROM2[4688]<=26'd11221774; ROM3[4688]<=26'd9750824; ROM4[4688]<=26'd23470555;
ROM1[4689]<=26'd1989871; ROM2[4689]<=26'd11230125; ROM3[4689]<=26'd9755157; ROM4[4689]<=26'd23475650;
ROM1[4690]<=26'd2005321; ROM2[4690]<=26'd11234465; ROM3[4690]<=26'd9750199; ROM4[4690]<=26'd23475675;
ROM1[4691]<=26'd2014581; ROM2[4691]<=26'd11236833; ROM3[4691]<=26'd9746368; ROM4[4691]<=26'd23476716;
ROM1[4692]<=26'd2007275; ROM2[4692]<=26'd11232409; ROM3[4692]<=26'd9744563; ROM4[4692]<=26'd23473933;
ROM1[4693]<=26'd1990276; ROM2[4693]<=26'd11224057; ROM3[4693]<=26'd9738457; ROM4[4693]<=26'd23466453;
ROM1[4694]<=26'd1983550; ROM2[4694]<=26'd11223644; ROM3[4694]<=26'd9741450; ROM4[4694]<=26'd23466696;
ROM1[4695]<=26'd1981303; ROM2[4695]<=26'd11226284; ROM3[4695]<=26'd9747342; ROM4[4695]<=26'd23469415;
ROM1[4696]<=26'd1982989; ROM2[4696]<=26'd11231153; ROM3[4696]<=26'd9750916; ROM4[4696]<=26'd23472524;
ROM1[4697]<=26'd1989917; ROM2[4697]<=26'd11234526; ROM3[4697]<=26'd9750032; ROM4[4697]<=26'd23473523;
ROM1[4698]<=26'd1998805; ROM2[4698]<=26'd11232855; ROM3[4698]<=26'd9743372; ROM4[4698]<=26'd23470046;
ROM1[4699]<=26'd2007394; ROM2[4699]<=26'd11233878; ROM3[4699]<=26'd9737632; ROM4[4699]<=26'd23468799;
ROM1[4700]<=26'd2007718; ROM2[4700]<=26'd11235674; ROM3[4700]<=26'd9739912; ROM4[4700]<=26'd23471120;
ROM1[4701]<=26'd2002206; ROM2[4701]<=26'd11235467; ROM3[4701]<=26'd9744916; ROM4[4701]<=26'd23472504;
ROM1[4702]<=26'd1995481; ROM2[4702]<=26'd11234791; ROM3[4702]<=26'd9748926; ROM4[4702]<=26'd23472787;
ROM1[4703]<=26'd1989957; ROM2[4703]<=26'd11235915; ROM3[4703]<=26'd9752685; ROM4[4703]<=26'd23474216;
ROM1[4704]<=26'd1983471; ROM2[4704]<=26'd11234030; ROM3[4704]<=26'd9755261; ROM4[4704]<=26'd23473464;
ROM1[4705]<=26'd1981658; ROM2[4705]<=26'd11228902; ROM3[4705]<=26'd9754712; ROM4[4705]<=26'd23471025;
ROM1[4706]<=26'd1987392; ROM2[4706]<=26'd11228399; ROM3[4706]<=26'd9749447; ROM4[4706]<=26'd23468873;
ROM1[4707]<=26'd1996357; ROM2[4707]<=26'd11228655; ROM3[4707]<=26'd9741725; ROM4[4707]<=26'd23465991;
ROM1[4708]<=26'd1998351; ROM2[4708]<=26'd11228351; ROM3[4708]<=26'd9740978; ROM4[4708]<=26'd23466266;
ROM1[4709]<=26'd1995111; ROM2[4709]<=26'd11229451; ROM3[4709]<=26'd9745058; ROM4[4709]<=26'd23467694;
ROM1[4710]<=26'd1987910; ROM2[4710]<=26'd11227568; ROM3[4710]<=26'd9749475; ROM4[4710]<=26'd23468297;
ROM1[4711]<=26'd1987020; ROM2[4711]<=26'd11228498; ROM3[4711]<=26'd9757122; ROM4[4711]<=26'd23472131;
ROM1[4712]<=26'd1987315; ROM2[4712]<=26'd11233224; ROM3[4712]<=26'd9765879; ROM4[4712]<=26'd23478549;
ROM1[4713]<=26'd1977504; ROM2[4713]<=26'd11226986; ROM3[4713]<=26'd9760057; ROM4[4713]<=26'd23472205;
ROM1[4714]<=26'd1976032; ROM2[4714]<=26'd11219062; ROM3[4714]<=26'd9750667; ROM4[4714]<=26'd23465482;
ROM1[4715]<=26'd1989414; ROM2[4715]<=26'd11220443; ROM3[4715]<=26'd9746073; ROM4[4715]<=26'd23465506;
ROM1[4716]<=26'd1998046; ROM2[4716]<=26'd11220698; ROM3[4716]<=26'd9743239; ROM4[4716]<=26'd23466222;
ROM1[4717]<=26'd2004482; ROM2[4717]<=26'd11228661; ROM3[4717]<=26'd9752985; ROM4[4717]<=26'd23475240;
ROM1[4718]<=26'd2006666; ROM2[4718]<=26'd11239063; ROM3[4718]<=26'd9764332; ROM4[4718]<=26'd23483041;
ROM1[4719]<=26'd1994126; ROM2[4719]<=26'd11232452; ROM3[4719]<=26'd9759418; ROM4[4719]<=26'd23476617;
ROM1[4720]<=26'd1979710; ROM2[4720]<=26'd11224908; ROM3[4720]<=26'd9752986; ROM4[4720]<=26'd23468123;
ROM1[4721]<=26'd1978955; ROM2[4721]<=26'd11227037; ROM3[4721]<=26'd9755076; ROM4[4721]<=26'd23470011;
ROM1[4722]<=26'd1982813; ROM2[4722]<=26'd11227619; ROM3[4722]<=26'd9752862; ROM4[4722]<=26'd23472212;
ROM1[4723]<=26'd1992394; ROM2[4723]<=26'd11225849; ROM3[4723]<=26'd9747460; ROM4[4723]<=26'd23471365;
ROM1[4724]<=26'd2002413; ROM2[4724]<=26'd11226052; ROM3[4724]<=26'd9739863; ROM4[4724]<=26'd23468656;
ROM1[4725]<=26'd1998257; ROM2[4725]<=26'd11227367; ROM3[4725]<=26'd9739835; ROM4[4725]<=26'd23470392;
ROM1[4726]<=26'd1994583; ROM2[4726]<=26'd11230722; ROM3[4726]<=26'd9746552; ROM4[4726]<=26'd23474701;
ROM1[4727]<=26'd1991947; ROM2[4727]<=26'd11233901; ROM3[4727]<=26'd9753258; ROM4[4727]<=26'd23477352;
ROM1[4728]<=26'd1982351; ROM2[4728]<=26'd11229093; ROM3[4728]<=26'd9753398; ROM4[4728]<=26'd23475557;
ROM1[4729]<=26'd1977773; ROM2[4729]<=26'd11223916; ROM3[4729]<=26'd9751112; ROM4[4729]<=26'd23470755;
ROM1[4730]<=26'd1982589; ROM2[4730]<=26'd11221968; ROM3[4730]<=26'd9750012; ROM4[4730]<=26'd23468909;
ROM1[4731]<=26'd1996231; ROM2[4731]<=26'd11225240; ROM3[4731]<=26'd9750886; ROM4[4731]<=26'd23472803;
ROM1[4732]<=26'd2007847; ROM2[4732]<=26'd11225928; ROM3[4732]<=26'd9748107; ROM4[4732]<=26'd23474219;
ROM1[4733]<=26'd2006571; ROM2[4733]<=26'd11224044; ROM3[4733]<=26'd9746969; ROM4[4733]<=26'd23472746;
ROM1[4734]<=26'd1998788; ROM2[4734]<=26'd11222433; ROM3[4734]<=26'd9749230; ROM4[4734]<=26'd23471888;
ROM1[4735]<=26'd1987962; ROM2[4735]<=26'd11220002; ROM3[4735]<=26'd9748509; ROM4[4735]<=26'd23469741;
ROM1[4736]<=26'd1990259; ROM2[4736]<=26'd11226921; ROM3[4736]<=26'd9757576; ROM4[4736]<=26'd23477119;
ROM1[4737]<=26'd1992645; ROM2[4737]<=26'd11234002; ROM3[4737]<=26'd9767186; ROM4[4737]<=26'd23484738;
ROM1[4738]<=26'd1987512; ROM2[4738]<=26'd11232571; ROM3[4738]<=26'd9763345; ROM4[4738]<=26'd23480775;
ROM1[4739]<=26'd1986629; ROM2[4739]<=26'd11227338; ROM3[4739]<=26'd9753787; ROM4[4739]<=26'd23472949;
ROM1[4740]<=26'd1999489; ROM2[4740]<=26'd11228948; ROM3[4740]<=26'd9745335; ROM4[4740]<=26'd23471020;
ROM1[4741]<=26'd2007828; ROM2[4741]<=26'd11230918; ROM3[4741]<=26'd9740559; ROM4[4741]<=26'd23470909;
ROM1[4742]<=26'd2005261; ROM2[4742]<=26'd11233021; ROM3[4742]<=26'd9743616; ROM4[4742]<=26'd23473400;
ROM1[4743]<=26'd2002203; ROM2[4743]<=26'd11236345; ROM3[4743]<=26'd9752216; ROM4[4743]<=26'd23478106;
ROM1[4744]<=26'd1994806; ROM2[4744]<=26'd11234708; ROM3[4744]<=26'd9757105; ROM4[4744]<=26'd23478013;
ROM1[4745]<=26'd1982984; ROM2[4745]<=26'd11229824; ROM3[4745]<=26'd9755722; ROM4[4745]<=26'd23475056;
ROM1[4746]<=26'd1976618; ROM2[4746]<=26'd11225864; ROM3[4746]<=26'd9754830; ROM4[4746]<=26'd23472706;
ROM1[4747]<=26'd1979867; ROM2[4747]<=26'd11226590; ROM3[4747]<=26'd9751623; ROM4[4747]<=26'd23470469;
ROM1[4748]<=26'd1991324; ROM2[4748]<=26'd11228764; ROM3[4748]<=26'd9746341; ROM4[4748]<=26'd23469829;
ROM1[4749]<=26'd2000344; ROM2[4749]<=26'd11227287; ROM3[4749]<=26'd9738848; ROM4[4749]<=26'd23466566;
ROM1[4750]<=26'd1993959; ROM2[4750]<=26'd11221919; ROM3[4750]<=26'd9733336; ROM4[4750]<=26'd23460614;
ROM1[4751]<=26'd1986221; ROM2[4751]<=26'd11221277; ROM3[4751]<=26'd9735253; ROM4[4751]<=26'd23461426;
ROM1[4752]<=26'd1983576; ROM2[4752]<=26'd11223383; ROM3[4752]<=26'd9739337; ROM4[4752]<=26'd23463376;
ROM1[4753]<=26'd1981751; ROM2[4753]<=26'd11226594; ROM3[4753]<=26'd9744501; ROM4[4753]<=26'd23465024;
ROM1[4754]<=26'd1978208; ROM2[4754]<=26'd11228775; ROM3[4754]<=26'd9747920; ROM4[4754]<=26'd23467640;
ROM1[4755]<=26'd1971654; ROM2[4755]<=26'd11221678; ROM3[4755]<=26'd9740539; ROM4[4755]<=26'd23459670;
ROM1[4756]<=26'd1969979; ROM2[4756]<=26'd11213322; ROM3[4756]<=26'd9729338; ROM4[4756]<=26'd23449091;
ROM1[4757]<=26'd1980158; ROM2[4757]<=26'd11212205; ROM3[4757]<=26'd9721638; ROM4[4757]<=26'd23446637;
ROM1[4758]<=26'd1983288; ROM2[4758]<=26'd11213737; ROM3[4758]<=26'd9720819; ROM4[4758]<=26'd23447352;
ROM1[4759]<=26'd1980744; ROM2[4759]<=26'd11216667; ROM3[4759]<=26'd9724764; ROM4[4759]<=26'd23451314;
ROM1[4760]<=26'd1977575; ROM2[4760]<=26'd11219175; ROM3[4760]<=26'd9731517; ROM4[4760]<=26'd23455221;
ROM1[4761]<=26'd1972860; ROM2[4761]<=26'd11218074; ROM3[4761]<=26'd9734787; ROM4[4761]<=26'd23455558;
ROM1[4762]<=26'd1967023; ROM2[4762]<=26'd11214864; ROM3[4762]<=26'd9737508; ROM4[4762]<=26'd23455828;
ROM1[4763]<=26'd1970287; ROM2[4763]<=26'd11215621; ROM3[4763]<=26'd9744031; ROM4[4763]<=26'd23459987;
ROM1[4764]<=26'd1977051; ROM2[4764]<=26'd11216991; ROM3[4764]<=26'd9742594; ROM4[4764]<=26'd23461147;
ROM1[4765]<=26'd1992196; ROM2[4765]<=26'd11220972; ROM3[4765]<=26'd9739962; ROM4[4765]<=26'd23464509;
ROM1[4766]<=26'd2003123; ROM2[4766]<=26'd11225275; ROM3[4766]<=26'd9739808; ROM4[4766]<=26'd23467903;
ROM1[4767]<=26'd1998619; ROM2[4767]<=26'd11225529; ROM3[4767]<=26'd9741019; ROM4[4767]<=26'd23467896;
ROM1[4768]<=26'd1991296; ROM2[4768]<=26'd11223349; ROM3[4768]<=26'd9745048; ROM4[4768]<=26'd23468098;
ROM1[4769]<=26'd1984071; ROM2[4769]<=26'd11221343; ROM3[4769]<=26'd9747159; ROM4[4769]<=26'd23466555;
ROM1[4770]<=26'd1976830; ROM2[4770]<=26'd11219540; ROM3[4770]<=26'd9748761; ROM4[4770]<=26'd23465128;
ROM1[4771]<=26'd1976912; ROM2[4771]<=26'd11221614; ROM3[4771]<=26'd9752155; ROM4[4771]<=26'd23466536;
ROM1[4772]<=26'd1990278; ROM2[4772]<=26'd11230885; ROM3[4772]<=26'd9757407; ROM4[4772]<=26'd23475307;
ROM1[4773]<=26'd2002950; ROM2[4773]<=26'd11233040; ROM3[4773]<=26'd9754749; ROM4[4773]<=26'd23478512;
ROM1[4774]<=26'd2006321; ROM2[4774]<=26'd11227042; ROM3[4774]<=26'd9743717; ROM4[4774]<=26'd23472072;
ROM1[4775]<=26'd1998226; ROM2[4775]<=26'd11221697; ROM3[4775]<=26'd9737595; ROM4[4775]<=26'd23466911;
ROM1[4776]<=26'd1988318; ROM2[4776]<=26'd11219343; ROM3[4776]<=26'd9739040; ROM4[4776]<=26'd23462987;
ROM1[4777]<=26'd1984347; ROM2[4777]<=26'd11219490; ROM3[4777]<=26'd9743992; ROM4[4777]<=26'd23462363;
ROM1[4778]<=26'd1983341; ROM2[4778]<=26'd11223295; ROM3[4778]<=26'd9747450; ROM4[4778]<=26'd23464995;
ROM1[4779]<=26'd1978489; ROM2[4779]<=26'd11223226; ROM3[4779]<=26'd9749271; ROM4[4779]<=26'd23465499;
ROM1[4780]<=26'd1976689; ROM2[4780]<=26'd11219656; ROM3[4780]<=26'd9746335; ROM4[4780]<=26'd23463616;
ROM1[4781]<=26'd1982916; ROM2[4781]<=26'd11219363; ROM3[4781]<=26'd9739615; ROM4[4781]<=26'd23461515;
ROM1[4782]<=26'd1996644; ROM2[4782]<=26'd11221624; ROM3[4782]<=26'd9736525; ROM4[4782]<=26'd23462555;
ROM1[4783]<=26'd2001185; ROM2[4783]<=26'd11224184; ROM3[4783]<=26'd9738118; ROM4[4783]<=26'd23464192;
ROM1[4784]<=26'd1994647; ROM2[4784]<=26'd11224730; ROM3[4784]<=26'd9739490; ROM4[4784]<=26'd23463808;
ROM1[4785]<=26'd1986969; ROM2[4785]<=26'd11223874; ROM3[4785]<=26'd9745048; ROM4[4785]<=26'd23465112;
ROM1[4786]<=26'd1983620; ROM2[4786]<=26'd11226472; ROM3[4786]<=26'd9751595; ROM4[4786]<=26'd23467453;
ROM1[4787]<=26'd1980026; ROM2[4787]<=26'd11226169; ROM3[4787]<=26'd9755153; ROM4[4787]<=26'd23469723;
ROM1[4788]<=26'd1980668; ROM2[4788]<=26'd11226220; ROM3[4788]<=26'd9755841; ROM4[4788]<=26'd23470160;
ROM1[4789]<=26'd1987304; ROM2[4789]<=26'd11227524; ROM3[4789]<=26'd9752401; ROM4[4789]<=26'd23469539;
ROM1[4790]<=26'd2002534; ROM2[4790]<=26'd11229489; ROM3[4790]<=26'd9750275; ROM4[4790]<=26'd23470866;
ROM1[4791]<=26'd2010174; ROM2[4791]<=26'd11230032; ROM3[4791]<=26'd9746143; ROM4[4791]<=26'd23468551;
ROM1[4792]<=26'd2002324; ROM2[4792]<=26'd11225570; ROM3[4792]<=26'd9743586; ROM4[4792]<=26'd23466172;
ROM1[4793]<=26'd2003258; ROM2[4793]<=26'd11233240; ROM3[4793]<=26'd9755546; ROM4[4793]<=26'd23475304;
ROM1[4794]<=26'd2002770; ROM2[4794]<=26'd11237732; ROM3[4794]<=26'd9762079; ROM4[4794]<=26'd23479103;
ROM1[4795]<=26'd1986227; ROM2[4795]<=26'd11224458; ROM3[4795]<=26'd9752189; ROM4[4795]<=26'd23468329;
ROM1[4796]<=26'd1971753; ROM2[4796]<=26'd11213661; ROM3[4796]<=26'd9742329; ROM4[4796]<=26'd23458118;
ROM1[4797]<=26'd1971858; ROM2[4797]<=26'd11210721; ROM3[4797]<=26'd9737815; ROM4[4797]<=26'd23454253;
ROM1[4798]<=26'd1984005; ROM2[4798]<=26'd11211895; ROM3[4798]<=26'd9736084; ROM4[4798]<=26'd23455848;
ROM1[4799]<=26'd2003087; ROM2[4799]<=26'd11223096; ROM3[4799]<=26'd9739554; ROM4[4799]<=26'd23464985;
ROM1[4800]<=26'd2007882; ROM2[4800]<=26'd11230512; ROM3[4800]<=26'd9745892; ROM4[4800]<=26'd23471520;
ROM1[4801]<=26'd1998942; ROM2[4801]<=26'd11227468; ROM3[4801]<=26'd9747472; ROM4[4801]<=26'd23469385;
ROM1[4802]<=26'd1992492; ROM2[4802]<=26'd11227366; ROM3[4802]<=26'd9749926; ROM4[4802]<=26'd23470224;
ROM1[4803]<=26'd1990424; ROM2[4803]<=26'd11229543; ROM3[4803]<=26'd9756639; ROM4[4803]<=26'd23475554;
ROM1[4804]<=26'd1987096; ROM2[4804]<=26'd11229143; ROM3[4804]<=26'd9761297; ROM4[4804]<=26'd23477535;
ROM1[4805]<=26'd1986166; ROM2[4805]<=26'd11226131; ROM3[4805]<=26'd9758527; ROM4[4805]<=26'd23474033;
ROM1[4806]<=26'd1989480; ROM2[4806]<=26'd11220664; ROM3[4806]<=26'd9747469; ROM4[4806]<=26'd23466753;
ROM1[4807]<=26'd1998837; ROM2[4807]<=26'd11218694; ROM3[4807]<=26'd9738592; ROM4[4807]<=26'd23463886;
ROM1[4808]<=26'd2004575; ROM2[4808]<=26'd11221869; ROM3[4808]<=26'd9740426; ROM4[4808]<=26'd23466861;
ROM1[4809]<=26'd2002930; ROM2[4809]<=26'd11224968; ROM3[4809]<=26'd9744429; ROM4[4809]<=26'd23471469;
ROM1[4810]<=26'd2000840; ROM2[4810]<=26'd11229240; ROM3[4810]<=26'd9753326; ROM4[4810]<=26'd23477567;
ROM1[4811]<=26'd2001278; ROM2[4811]<=26'd11233357; ROM3[4811]<=26'd9762566; ROM4[4811]<=26'd23482715;
ROM1[4812]<=26'd1990774; ROM2[4812]<=26'd11227480; ROM3[4812]<=26'd9759296; ROM4[4812]<=26'd23477406;
ROM1[4813]<=26'd1977283; ROM2[4813]<=26'd11216590; ROM3[4813]<=26'd9750168; ROM4[4813]<=26'd23465573;
ROM1[4814]<=26'd1977937; ROM2[4814]<=26'd11211784; ROM3[4814]<=26'd9742985; ROM4[4814]<=26'd23460946;
ROM1[4815]<=26'd1989187; ROM2[4815]<=26'd11211035; ROM3[4815]<=26'd9736464; ROM4[4815]<=26'd23458741;
ROM1[4816]<=26'd1996942; ROM2[4816]<=26'd11213225; ROM3[4816]<=26'd9735071; ROM4[4816]<=26'd23460304;
ROM1[4817]<=26'd1993879; ROM2[4817]<=26'd11214012; ROM3[4817]<=26'd9736405; ROM4[4817]<=26'd23463295;
ROM1[4818]<=26'd1986891; ROM2[4818]<=26'd11213206; ROM3[4818]<=26'd9740647; ROM4[4818]<=26'd23464874;
ROM1[4819]<=26'd1982002; ROM2[4819]<=26'd11213990; ROM3[4819]<=26'd9745722; ROM4[4819]<=26'd23466046;
ROM1[4820]<=26'd1980931; ROM2[4820]<=26'd11217294; ROM3[4820]<=26'd9754199; ROM4[4820]<=26'd23470507;
ROM1[4821]<=26'd1983947; ROM2[4821]<=26'd11220857; ROM3[4821]<=26'd9762815; ROM4[4821]<=26'd23477416;
ROM1[4822]<=26'd1989810; ROM2[4822]<=26'd11225816; ROM3[4822]<=26'd9763303; ROM4[4822]<=26'd23478952;
ROM1[4823]<=26'd1997027; ROM2[4823]<=26'd11224271; ROM3[4823]<=26'd9756960; ROM4[4823]<=26'd23474419;
ROM1[4824]<=26'd2003263; ROM2[4824]<=26'd11220231; ROM3[4824]<=26'd9748838; ROM4[4824]<=26'd23470063;
ROM1[4825]<=26'd2001747; ROM2[4825]<=26'd11221654; ROM3[4825]<=26'd9747764; ROM4[4825]<=26'd23469892;
ROM1[4826]<=26'd1993047; ROM2[4826]<=26'd11218964; ROM3[4826]<=26'd9749233; ROM4[4826]<=26'd23468307;
ROM1[4827]<=26'd1986084; ROM2[4827]<=26'd11217737; ROM3[4827]<=26'd9751629; ROM4[4827]<=26'd23467666;
ROM1[4828]<=26'd1982822; ROM2[4828]<=26'd11220201; ROM3[4828]<=26'd9756254; ROM4[4828]<=26'd23470560;
ROM1[4829]<=26'd1982682; ROM2[4829]<=26'd11223367; ROM3[4829]<=26'd9764467; ROM4[4829]<=26'd23474364;
ROM1[4830]<=26'd1981776; ROM2[4830]<=26'd11219816; ROM3[4830]<=26'd9759722; ROM4[4830]<=26'd23470768;
ROM1[4831]<=26'd1984230; ROM2[4831]<=26'd11213826; ROM3[4831]<=26'd9749565; ROM4[4831]<=26'd23464178;
ROM1[4832]<=26'd1998945; ROM2[4832]<=26'd11216363; ROM3[4832]<=26'd9747120; ROM4[4832]<=26'd23466395;
ROM1[4833]<=26'd2002060; ROM2[4833]<=26'd11217426; ROM3[4833]<=26'd9745293; ROM4[4833]<=26'd23468089;
ROM1[4834]<=26'd1994615; ROM2[4834]<=26'd11216200; ROM3[4834]<=26'd9749267; ROM4[4834]<=26'd23468288;
ROM1[4835]<=26'd1988951; ROM2[4835]<=26'd11216011; ROM3[4835]<=26'd9754944; ROM4[4835]<=26'd23470037;
ROM1[4836]<=26'd1990497; ROM2[4836]<=26'd11220963; ROM3[4836]<=26'd9760591; ROM4[4836]<=26'd23473448;
ROM1[4837]<=26'd1997989; ROM2[4837]<=26'd11234134; ROM3[4837]<=26'd9775466; ROM4[4837]<=26'd23485589;
ROM1[4838]<=26'd1998332; ROM2[4838]<=26'd11233912; ROM3[4838]<=26'd9776142; ROM4[4838]<=26'd23485363;
ROM1[4839]<=26'd1989576; ROM2[4839]<=26'd11220089; ROM3[4839]<=26'd9758967; ROM4[4839]<=26'd23470254;
ROM1[4840]<=26'd1996313; ROM2[4840]<=26'd11215924; ROM3[4840]<=26'd9750156; ROM4[4840]<=26'd23465968;
ROM1[4841]<=26'd1994715; ROM2[4841]<=26'd11209599; ROM3[4841]<=26'd9738405; ROM4[4841]<=26'd23458403;
ROM1[4842]<=26'd1991094; ROM2[4842]<=26'd11209277; ROM3[4842]<=26'd9739357; ROM4[4842]<=26'd23459894;
ROM1[4843]<=26'd1994655; ROM2[4843]<=26'd11221402; ROM3[4843]<=26'd9754255; ROM4[4843]<=26'd23472736;
ROM1[4844]<=26'd1990412; ROM2[4844]<=26'd11224534; ROM3[4844]<=26'd9759767; ROM4[4844]<=26'd23474690;
ROM1[4845]<=26'd1978704; ROM2[4845]<=26'd11215188; ROM3[4845]<=26'd9755371; ROM4[4845]<=26'd23467443;
ROM1[4846]<=26'd1971708; ROM2[4846]<=26'd11211739; ROM3[4846]<=26'd9753206; ROM4[4846]<=26'd23464587;
ROM1[4847]<=26'd1980128; ROM2[4847]<=26'd11217265; ROM3[4847]<=26'd9756152; ROM4[4847]<=26'd23469224;
ROM1[4848]<=26'd1991974; ROM2[4848]<=26'd11218518; ROM3[4848]<=26'd9750221; ROM4[4848]<=26'd23468388;
ROM1[4849]<=26'd2002718; ROM2[4849]<=26'd11218889; ROM3[4849]<=26'd9744658; ROM4[4849]<=26'd23467728;
ROM1[4850]<=26'd2003037; ROM2[4850]<=26'd11221666; ROM3[4850]<=26'd9745597; ROM4[4850]<=26'd23470746;
ROM1[4851]<=26'd1996990; ROM2[4851]<=26'd11222755; ROM3[4851]<=26'd9750091; ROM4[4851]<=26'd23472846;
ROM1[4852]<=26'd1990127; ROM2[4852]<=26'd11221330; ROM3[4852]<=26'd9754386; ROM4[4852]<=26'd23474178;
ROM1[4853]<=26'd1980635; ROM2[4853]<=26'd11218485; ROM3[4853]<=26'd9753582; ROM4[4853]<=26'd23471085;
ROM1[4854]<=26'd1964455; ROM2[4854]<=26'd11210107; ROM3[4854]<=26'd9746957; ROM4[4854]<=26'd23461387;
ROM1[4855]<=26'd1965096; ROM2[4855]<=26'd11208427; ROM3[4855]<=26'd9742607; ROM4[4855]<=26'd23457744;
ROM1[4856]<=26'd1974712; ROM2[4856]<=26'd11208525; ROM3[4856]<=26'd9738682; ROM4[4856]<=26'd23456949;
ROM1[4857]<=26'd1986357; ROM2[4857]<=26'd11211390; ROM3[4857]<=26'd9735796; ROM4[4857]<=26'd23459179;
ROM1[4858]<=26'd1995833; ROM2[4858]<=26'd11216949; ROM3[4858]<=26'd9739889; ROM4[4858]<=26'd23463912;
ROM1[4859]<=26'd1992567; ROM2[4859]<=26'd11217323; ROM3[4859]<=26'd9744200; ROM4[4859]<=26'd23466043;
ROM1[4860]<=26'd1983002; ROM2[4860]<=26'd11217317; ROM3[4860]<=26'd9747487; ROM4[4860]<=26'd23464941;
ROM1[4861]<=26'd1975095; ROM2[4861]<=26'd11213397; ROM3[4861]<=26'd9745647; ROM4[4861]<=26'd23459467;
ROM1[4862]<=26'd1973740; ROM2[4862]<=26'd11216038; ROM3[4862]<=26'd9751051; ROM4[4862]<=26'd23464840;
ROM1[4863]<=26'd1973037; ROM2[4863]<=26'd11217643; ROM3[4863]<=26'd9752143; ROM4[4863]<=26'd23466797;
ROM1[4864]<=26'd1975515; ROM2[4864]<=26'd11213378; ROM3[4864]<=26'd9744051; ROM4[4864]<=26'd23461062;
ROM1[4865]<=26'd1987485; ROM2[4865]<=26'd11214148; ROM3[4865]<=26'd9739232; ROM4[4865]<=26'd23460877;
ROM1[4866]<=26'd1992587; ROM2[4866]<=26'd11213341; ROM3[4866]<=26'd9734491; ROM4[4866]<=26'd23458868;
ROM1[4867]<=26'd1988075; ROM2[4867]<=26'd11211093; ROM3[4867]<=26'd9734810; ROM4[4867]<=26'd23459512;
ROM1[4868]<=26'd1979527; ROM2[4868]<=26'd11209584; ROM3[4868]<=26'd9736862; ROM4[4868]<=26'd23459281;
ROM1[4869]<=26'd1974161; ROM2[4869]<=26'd11208417; ROM3[4869]<=26'd9738284; ROM4[4869]<=26'd23457599;
ROM1[4870]<=26'd1969765; ROM2[4870]<=26'd11207576; ROM3[4870]<=26'd9742943; ROM4[4870]<=26'd23457614;
ROM1[4871]<=26'd1966468; ROM2[4871]<=26'd11207319; ROM3[4871]<=26'd9745817; ROM4[4871]<=26'd23457552;
ROM1[4872]<=26'd1971121; ROM2[4872]<=26'd11210765; ROM3[4872]<=26'd9745546; ROM4[4872]<=26'd23459613;
ROM1[4873]<=26'd1982666; ROM2[4873]<=26'd11213216; ROM3[4873]<=26'd9743069; ROM4[4873]<=26'd23460186;
ROM1[4874]<=26'd1994674; ROM2[4874]<=26'd11214311; ROM3[4874]<=26'd9740883; ROM4[4874]<=26'd23461523;
ROM1[4875]<=26'd1996027; ROM2[4875]<=26'd11216689; ROM3[4875]<=26'd9743157; ROM4[4875]<=26'd23462996;
ROM1[4876]<=26'd1990372; ROM2[4876]<=26'd11214352; ROM3[4876]<=26'd9746577; ROM4[4876]<=26'd23463592;
ROM1[4877]<=26'd1986889; ROM2[4877]<=26'd11215400; ROM3[4877]<=26'd9752262; ROM4[4877]<=26'd23466954;
ROM1[4878]<=26'd1983957; ROM2[4878]<=26'd11219392; ROM3[4878]<=26'd9757897; ROM4[4878]<=26'd23470099;
ROM1[4879]<=26'd1980790; ROM2[4879]<=26'd11221671; ROM3[4879]<=26'd9762381; ROM4[4879]<=26'd23473136;
ROM1[4880]<=26'd1980007; ROM2[4880]<=26'd11219725; ROM3[4880]<=26'd9760000; ROM4[4880]<=26'd23472126;
ROM1[4881]<=26'd1986139; ROM2[4881]<=26'd11215851; ROM3[4881]<=26'd9752381; ROM4[4881]<=26'd23468843;
ROM1[4882]<=26'd1995848; ROM2[4882]<=26'd11213710; ROM3[4882]<=26'd9743012; ROM4[4882]<=26'd23464488;
ROM1[4883]<=26'd1992700; ROM2[4883]<=26'd11209228; ROM3[4883]<=26'd9737702; ROM4[4883]<=26'd23459640;
ROM1[4884]<=26'd1988316; ROM2[4884]<=26'd11211944; ROM3[4884]<=26'd9742234; ROM4[4884]<=26'd23461664;
ROM1[4885]<=26'd1983760; ROM2[4885]<=26'd11214794; ROM3[4885]<=26'd9748052; ROM4[4885]<=26'd23463902;
ROM1[4886]<=26'd1974947; ROM2[4886]<=26'd11210851; ROM3[4886]<=26'd9747604; ROM4[4886]<=26'd23461410;
ROM1[4887]<=26'd1965343; ROM2[4887]<=26'd11206096; ROM3[4887]<=26'd9747209; ROM4[4887]<=26'd23459160;
ROM1[4888]<=26'd1962365; ROM2[4888]<=26'd11203429; ROM3[4888]<=26'd9746202; ROM4[4888]<=26'd23456888;
ROM1[4889]<=26'd1969264; ROM2[4889]<=26'd11205144; ROM3[4889]<=26'd9744172; ROM4[4889]<=26'd23456444;
ROM1[4890]<=26'd1984967; ROM2[4890]<=26'd11208422; ROM3[4890]<=26'd9743162; ROM4[4890]<=26'd23459688;
ROM1[4891]<=26'd1993660; ROM2[4891]<=26'd11211688; ROM3[4891]<=26'd9742071; ROM4[4891]<=26'd23463434;
ROM1[4892]<=26'd1994919; ROM2[4892]<=26'd11217781; ROM3[4892]<=26'd9748711; ROM4[4892]<=26'd23469726;
ROM1[4893]<=26'd1994322; ROM2[4893]<=26'd11221529; ROM3[4893]<=26'd9759197; ROM4[4893]<=26'd23476135;
ROM1[4894]<=26'd1982179; ROM2[4894]<=26'd11215414; ROM3[4894]<=26'd9757569; ROM4[4894]<=26'd23470738;
ROM1[4895]<=26'd1971645; ROM2[4895]<=26'd11209030; ROM3[4895]<=26'd9755500; ROM4[4895]<=26'd23464636;
ROM1[4896]<=26'd1966794; ROM2[4896]<=26'd11204941; ROM3[4896]<=26'd9753477; ROM4[4896]<=26'd23461413;
ROM1[4897]<=26'd1965355; ROM2[4897]<=26'd11201151; ROM3[4897]<=26'd9748410; ROM4[4897]<=26'd23457490;
ROM1[4898]<=26'd1984664; ROM2[4898]<=26'd11208525; ROM3[4898]<=26'd9752408; ROM4[4898]<=26'd23464663;
ROM1[4899]<=26'd1993832; ROM2[4899]<=26'd11208915; ROM3[4899]<=26'd9746436; ROM4[4899]<=26'd23463130;
ROM1[4900]<=26'd1981617; ROM2[4900]<=26'd11201127; ROM3[4900]<=26'd9740053; ROM4[4900]<=26'd23454922;
ROM1[4901]<=26'd1973091; ROM2[4901]<=26'd11200659; ROM3[4901]<=26'd9743285; ROM4[4901]<=26'd23456578;
ROM1[4902]<=26'd1967854; ROM2[4902]<=26'd11201801; ROM3[4902]<=26'd9746995; ROM4[4902]<=26'd23457989;
ROM1[4903]<=26'd1969256; ROM2[4903]<=26'd11206042; ROM3[4903]<=26'd9755369; ROM4[4903]<=26'd23463416;
ROM1[4904]<=26'd1970792; ROM2[4904]<=26'd11210420; ROM3[4904]<=26'd9760999; ROM4[4904]<=26'd23469544;
ROM1[4905]<=26'd1971531; ROM2[4905]<=26'd11209658; ROM3[4905]<=26'd9759055; ROM4[4905]<=26'd23466345;
ROM1[4906]<=26'd1979606; ROM2[4906]<=26'd11209696; ROM3[4906]<=26'd9753206; ROM4[4906]<=26'd23463466;
ROM1[4907]<=26'd1994406; ROM2[4907]<=26'd11211467; ROM3[4907]<=26'd9747744; ROM4[4907]<=26'd23464414;
ROM1[4908]<=26'd1996386; ROM2[4908]<=26'd11209813; ROM3[4908]<=26'd9745750; ROM4[4908]<=26'd23463662;
ROM1[4909]<=26'd1988530; ROM2[4909]<=26'd11208664; ROM3[4909]<=26'd9747472; ROM4[4909]<=26'd23463331;
ROM1[4910]<=26'd1982100; ROM2[4910]<=26'd11209768; ROM3[4910]<=26'd9752342; ROM4[4910]<=26'd23467200;
ROM1[4911]<=26'd1979115; ROM2[4911]<=26'd11212375; ROM3[4911]<=26'd9757906; ROM4[4911]<=26'd23470298;
ROM1[4912]<=26'd1974540; ROM2[4912]<=26'd11212734; ROM3[4912]<=26'd9761946; ROM4[4912]<=26'd23471183;
ROM1[4913]<=26'd1971007; ROM2[4913]<=26'd11209787; ROM3[4913]<=26'd9760664; ROM4[4913]<=26'd23470400;
ROM1[4914]<=26'd1974927; ROM2[4914]<=26'd11207996; ROM3[4914]<=26'd9756711; ROM4[4914]<=26'd23467178;
ROM1[4915]<=26'd1990693; ROM2[4915]<=26'd11212753; ROM3[4915]<=26'd9754299; ROM4[4915]<=26'd23469286;
ROM1[4916]<=26'd2004765; ROM2[4916]<=26'd11219031; ROM3[4916]<=26'd9755953; ROM4[4916]<=26'd23474589;
ROM1[4917]<=26'd2000462; ROM2[4917]<=26'd11218442; ROM3[4917]<=26'd9755653; ROM4[4917]<=26'd23473499;
ROM1[4918]<=26'd1986572; ROM2[4918]<=26'd11212846; ROM3[4918]<=26'd9753032; ROM4[4918]<=26'd23468229;
ROM1[4919]<=26'd1978284; ROM2[4919]<=26'd11210437; ROM3[4919]<=26'd9754120; ROM4[4919]<=26'd23466385;
ROM1[4920]<=26'd1971324; ROM2[4920]<=26'd11210735; ROM3[4920]<=26'd9755870; ROM4[4920]<=26'd23465885;
ROM1[4921]<=26'd1971198; ROM2[4921]<=26'd11211936; ROM3[4921]<=26'd9759144; ROM4[4921]<=26'd23467473;
ROM1[4922]<=26'd1976085; ROM2[4922]<=26'd11211576; ROM3[4922]<=26'd9755496; ROM4[4922]<=26'd23467203;
ROM1[4923]<=26'd1984133; ROM2[4923]<=26'd11208613; ROM3[4923]<=26'd9747132; ROM4[4923]<=26'd23462922;
ROM1[4924]<=26'd1994972; ROM2[4924]<=26'd11207483; ROM3[4924]<=26'd9742704; ROM4[4924]<=26'd23462798;
ROM1[4925]<=26'd1996277; ROM2[4925]<=26'd11210386; ROM3[4925]<=26'd9745664; ROM4[4925]<=26'd23468198;
ROM1[4926]<=26'd1996922; ROM2[4926]<=26'd11216878; ROM3[4926]<=26'd9758028; ROM4[4926]<=26'd23475696;
ROM1[4927]<=26'd1987085; ROM2[4927]<=26'd11212752; ROM3[4927]<=26'd9760136; ROM4[4927]<=26'd23473666;
ROM1[4928]<=26'd1971623; ROM2[4928]<=26'd11204151; ROM3[4928]<=26'd9754729; ROM4[4928]<=26'd23466924;
ROM1[4929]<=26'd1967594; ROM2[4929]<=26'd11205931; ROM3[4929]<=26'd9755290; ROM4[4929]<=26'd23465257;
ROM1[4930]<=26'd1969914; ROM2[4930]<=26'd11207747; ROM3[4930]<=26'd9751655; ROM4[4930]<=26'd23463417;
ROM1[4931]<=26'd1981378; ROM2[4931]<=26'd11211238; ROM3[4931]<=26'd9746417; ROM4[4931]<=26'd23463651;
ROM1[4932]<=26'd1997146; ROM2[4932]<=26'd11215537; ROM3[4932]<=26'd9743014; ROM4[4932]<=26'd23464171;
ROM1[4933]<=26'd2001264; ROM2[4933]<=26'd11215506; ROM3[4933]<=26'd9742280; ROM4[4933]<=26'd23464910;
ROM1[4934]<=26'd1991352; ROM2[4934]<=26'd11209721; ROM3[4934]<=26'd9739334; ROM4[4934]<=26'd23461792;
ROM1[4935]<=26'd1983367; ROM2[4935]<=26'd11208309; ROM3[4935]<=26'd9743487; ROM4[4935]<=26'd23460713;
ROM1[4936]<=26'd1984955; ROM2[4936]<=26'd11214990; ROM3[4936]<=26'd9753549; ROM4[4936]<=26'd23468546;
ROM1[4937]<=26'd1975604; ROM2[4937]<=26'd11211301; ROM3[4937]<=26'd9752483; ROM4[4937]<=26'd23465467;
ROM1[4938]<=26'd1969290; ROM2[4938]<=26'd11205888; ROM3[4938]<=26'd9746549; ROM4[4938]<=26'd23458301;
ROM1[4939]<=26'd1978515; ROM2[4939]<=26'd11208912; ROM3[4939]<=26'd9743974; ROM4[4939]<=26'd23459696;
ROM1[4940]<=26'd1990181; ROM2[4940]<=26'd11209336; ROM3[4940]<=26'd9736838; ROM4[4940]<=26'd23456757;
ROM1[4941]<=26'd1998412; ROM2[4941]<=26'd11210566; ROM3[4941]<=26'd9733461; ROM4[4941]<=26'd23457898;
ROM1[4942]<=26'd2004454; ROM2[4942]<=26'd11218444; ROM3[4942]<=26'd9743777; ROM4[4942]<=26'd23466652;
ROM1[4943]<=26'd1995480; ROM2[4943]<=26'd11216663; ROM3[4943]<=26'd9747375; ROM4[4943]<=26'd23466706;
ROM1[4944]<=26'd1986538; ROM2[4944]<=26'd11213471; ROM3[4944]<=26'd9746940; ROM4[4944]<=26'd23464050;
ROM1[4945]<=26'd1979710; ROM2[4945]<=26'd11211554; ROM3[4945]<=26'd9750974; ROM4[4945]<=26'd23463258;
ROM1[4946]<=26'd1975684; ROM2[4946]<=26'd11212145; ROM3[4946]<=26'd9753988; ROM4[4946]<=26'd23465569;
ROM1[4947]<=26'd1985306; ROM2[4947]<=26'd11218457; ROM3[4947]<=26'd9756621; ROM4[4947]<=26'd23470278;
ROM1[4948]<=26'd1995844; ROM2[4948]<=26'd11217718; ROM3[4948]<=26'd9751680; ROM4[4948]<=26'd23469267;
ROM1[4949]<=26'd2003956; ROM2[4949]<=26'd11217037; ROM3[4949]<=26'd9744010; ROM4[4949]<=26'd23466934;
ROM1[4950]<=26'd2000067; ROM2[4950]<=26'd11214868; ROM3[4950]<=26'd9743439; ROM4[4950]<=26'd23466179;
ROM1[4951]<=26'd1989197; ROM2[4951]<=26'd11208103; ROM3[4951]<=26'd9742814; ROM4[4951]<=26'd23462934;
ROM1[4952]<=26'd1983966; ROM2[4952]<=26'd11207324; ROM3[4952]<=26'd9747696; ROM4[4952]<=26'd23463733;
ROM1[4953]<=26'd1977753; ROM2[4953]<=26'd11206798; ROM3[4953]<=26'd9750313; ROM4[4953]<=26'd23463187;
ROM1[4954]<=26'd1973328; ROM2[4954]<=26'd11206515; ROM3[4954]<=26'd9750901; ROM4[4954]<=26'd23462104;
ROM1[4955]<=26'd1976331; ROM2[4955]<=26'd11209151; ROM3[4955]<=26'd9752422; ROM4[4955]<=26'd23463245;
ROM1[4956]<=26'd1988205; ROM2[4956]<=26'd11214187; ROM3[4956]<=26'd9752212; ROM4[4956]<=26'd23466204;
ROM1[4957]<=26'd1999874; ROM2[4957]<=26'd11215194; ROM3[4957]<=26'd9746599; ROM4[4957]<=26'd23466298;
ROM1[4958]<=26'd1993481; ROM2[4958]<=26'd11205974; ROM3[4958]<=26'd9735750; ROM4[4958]<=26'd23458379;
ROM1[4959]<=26'd1987261; ROM2[4959]<=26'd11206029; ROM3[4959]<=26'd9736980; ROM4[4959]<=26'd23458722;
ROM1[4960]<=26'd1980385; ROM2[4960]<=26'd11204502; ROM3[4960]<=26'd9739111; ROM4[4960]<=26'd23460035;
ROM1[4961]<=26'd1976497; ROM2[4961]<=26'd11203055; ROM3[4961]<=26'd9739758; ROM4[4961]<=26'd23460120;
ROM1[4962]<=26'd1976516; ROM2[4962]<=26'd11209395; ROM3[4962]<=26'd9747101; ROM4[4962]<=26'd23465203;
ROM1[4963]<=26'd1974588; ROM2[4963]<=26'd11209017; ROM3[4963]<=26'd9746660; ROM4[4963]<=26'd23464198;
ROM1[4964]<=26'd1979135; ROM2[4964]<=26'd11208069; ROM3[4964]<=26'd9741955; ROM4[4964]<=26'd23462534;
ROM1[4965]<=26'd1993686; ROM2[4965]<=26'd11211109; ROM3[4965]<=26'd9738018; ROM4[4965]<=26'd23464315;
ROM1[4966]<=26'd2000291; ROM2[4966]<=26'd11211436; ROM3[4966]<=26'd9735448; ROM4[4966]<=26'd23464834;
ROM1[4967]<=26'd1994415; ROM2[4967]<=26'd11207738; ROM3[4967]<=26'd9735081; ROM4[4967]<=26'd23462648;
ROM1[4968]<=26'd1986763; ROM2[4968]<=26'd11206237; ROM3[4968]<=26'd9737426; ROM4[4968]<=26'd23461079;
ROM1[4969]<=26'd1979855; ROM2[4969]<=26'd11205163; ROM3[4969]<=26'd9742225; ROM4[4969]<=26'd23462005;
ROM1[4970]<=26'd1974558; ROM2[4970]<=26'd11206197; ROM3[4970]<=26'd9747155; ROM4[4970]<=26'd23462579;
ROM1[4971]<=26'd1971619; ROM2[4971]<=26'd11206959; ROM3[4971]<=26'd9749149; ROM4[4971]<=26'd23463130;
ROM1[4972]<=26'd1974236; ROM2[4972]<=26'd11206229; ROM3[4972]<=26'd9744700; ROM4[4972]<=26'd23461121;
ROM1[4973]<=26'd1984031; ROM2[4973]<=26'd11207469; ROM3[4973]<=26'd9739919; ROM4[4973]<=26'd23459486;
ROM1[4974]<=26'd1994822; ROM2[4974]<=26'd11207801; ROM3[4974]<=26'd9737539; ROM4[4974]<=26'd23460315;
ROM1[4975]<=26'd1995887; ROM2[4975]<=26'd11209698; ROM3[4975]<=26'd9739313; ROM4[4975]<=26'd23463134;
ROM1[4976]<=26'd1991549; ROM2[4976]<=26'd11212676; ROM3[4976]<=26'd9745021; ROM4[4976]<=26'd23465977;
ROM1[4977]<=26'd1986661; ROM2[4977]<=26'd11211194; ROM3[4977]<=26'd9748880; ROM4[4977]<=26'd23465492;
ROM1[4978]<=26'd1978016; ROM2[4978]<=26'd11207873; ROM3[4978]<=26'd9747136; ROM4[4978]<=26'd23461723;
ROM1[4979]<=26'd1970296; ROM2[4979]<=26'd11204340; ROM3[4979]<=26'd9745297; ROM4[4979]<=26'd23458704;
ROM1[4980]<=26'd1972407; ROM2[4980]<=26'd11204538; ROM3[4980]<=26'd9746443; ROM4[4980]<=26'd23458930;
ROM1[4981]<=26'd1982832; ROM2[4981]<=26'd11207845; ROM3[4981]<=26'd9743790; ROM4[4981]<=26'd23460277;
ROM1[4982]<=26'd1995164; ROM2[4982]<=26'd11207650; ROM3[4982]<=26'd9737383; ROM4[4982]<=26'd23459249;
ROM1[4983]<=26'd1995518; ROM2[4983]<=26'd11206696; ROM3[4983]<=26'd9733307; ROM4[4983]<=26'd23456172;
ROM1[4984]<=26'd1989821; ROM2[4984]<=26'd11206459; ROM3[4984]<=26'd9734268; ROM4[4984]<=26'd23456843;
ROM1[4985]<=26'd1988697; ROM2[4985]<=26'd11210450; ROM3[4985]<=26'd9743663; ROM4[4985]<=26'd23463896;
ROM1[4986]<=26'd1990555; ROM2[4986]<=26'd11217475; ROM3[4986]<=26'd9753675; ROM4[4986]<=26'd23472442;
ROM1[4987]<=26'd1988635; ROM2[4987]<=26'd11220306; ROM3[4987]<=26'd9761495; ROM4[4987]<=26'd23477147;
ROM1[4988]<=26'd1988959; ROM2[4988]<=26'd11220425; ROM3[4988]<=26'd9762229; ROM4[4988]<=26'd23476004;
ROM1[4989]<=26'd1992870; ROM2[4989]<=26'd11218519; ROM3[4989]<=26'd9755209; ROM4[4989]<=26'd23472464;
ROM1[4990]<=26'd1994645; ROM2[4990]<=26'd11209979; ROM3[4990]<=26'd9741899; ROM4[4990]<=26'd23462787;
ROM1[4991]<=26'd1993805; ROM2[4991]<=26'd11203991; ROM3[4991]<=26'd9733684; ROM4[4991]<=26'd23455615;
ROM1[4992]<=26'd1985669; ROM2[4992]<=26'd11200195; ROM3[4992]<=26'd9732284; ROM4[4992]<=26'd23452685;
ROM1[4993]<=26'd1976669; ROM2[4993]<=26'd11199184; ROM3[4993]<=26'd9734725; ROM4[4993]<=26'd23451131;
ROM1[4994]<=26'd1978377; ROM2[4994]<=26'd11206734; ROM3[4994]<=26'd9743002; ROM4[4994]<=26'd23457568;
ROM1[4995]<=26'd1979543; ROM2[4995]<=26'd11212032; ROM3[4995]<=26'd9750196; ROM4[4995]<=26'd23463550;
ROM1[4996]<=26'd1982756; ROM2[4996]<=26'd11216832; ROM3[4996]<=26'd9757654; ROM4[4996]<=26'd23469387;
ROM1[4997]<=26'd1983279; ROM2[4997]<=26'd11212827; ROM3[4997]<=26'd9754406; ROM4[4997]<=26'd23466078;
ROM1[4998]<=26'd1984211; ROM2[4998]<=26'd11203447; ROM3[4998]<=26'd9741030; ROM4[4998]<=26'd23456595;
ROM1[4999]<=26'd1993447; ROM2[4999]<=26'd11204107; ROM3[4999]<=26'd9736244; ROM4[4999]<=26'd23456837;
ROM1[5000]<=26'd1991460; ROM2[5000]<=26'd11204434; ROM3[5000]<=26'd9736562; ROM4[5000]<=26'd23457195;
ROM1[5001]<=26'd1987124; ROM2[5001]<=26'd11205502; ROM3[5001]<=26'd9742683; ROM4[5001]<=26'd23459907;
ROM1[5002]<=26'd1989451; ROM2[5002]<=26'd11211882; ROM3[5002]<=26'd9754522; ROM4[5002]<=26'd23468111;
ROM1[5003]<=26'd1982627; ROM2[5003]<=26'd11211153; ROM3[5003]<=26'd9756281; ROM4[5003]<=26'd23468665;
ROM1[5004]<=26'd1973633; ROM2[5004]<=26'd11207118; ROM3[5004]<=26'd9755435; ROM4[5004]<=26'd23464994;
ROM1[5005]<=26'd1974860; ROM2[5005]<=26'd11209140; ROM3[5005]<=26'd9752838; ROM4[5005]<=26'd23463363;
ROM1[5006]<=26'd1987270; ROM2[5006]<=26'd11212828; ROM3[5006]<=26'd9750266; ROM4[5006]<=26'd23464465;
ROM1[5007]<=26'd1998680; ROM2[5007]<=26'd11212223; ROM3[5007]<=26'd9743358; ROM4[5007]<=26'd23461618;
ROM1[5008]<=26'd1996798; ROM2[5008]<=26'd11208270; ROM3[5008]<=26'd9738884; ROM4[5008]<=26'd23457926;
ROM1[5009]<=26'd1990483; ROM2[5009]<=26'd11206860; ROM3[5009]<=26'd9741287; ROM4[5009]<=26'd23459014;
ROM1[5010]<=26'd1981500; ROM2[5010]<=26'd11205414; ROM3[5010]<=26'd9744107; ROM4[5010]<=26'd23459041;
ROM1[5011]<=26'd1977492; ROM2[5011]<=26'd11207601; ROM3[5011]<=26'd9747924; ROM4[5011]<=26'd23459371;
ROM1[5012]<=26'd1973342; ROM2[5012]<=26'd11209664; ROM3[5012]<=26'd9750176; ROM4[5012]<=26'd23460912;
ROM1[5013]<=26'd1972671; ROM2[5013]<=26'd11206174; ROM3[5013]<=26'd9748953; ROM4[5013]<=26'd23459304;
ROM1[5014]<=26'd1982089; ROM2[5014]<=26'd11207677; ROM3[5014]<=26'd9747835; ROM4[5014]<=26'd23460822;
ROM1[5015]<=26'd1998573; ROM2[5015]<=26'd11211894; ROM3[5015]<=26'd9747088; ROM4[5015]<=26'd23465261;
ROM1[5016]<=26'd2006721; ROM2[5016]<=26'd11213762; ROM3[5016]<=26'd9746619; ROM4[5016]<=26'd23466637;
ROM1[5017]<=26'd2001833; ROM2[5017]<=26'd11214370; ROM3[5017]<=26'd9747450; ROM4[5017]<=26'd23465608;
ROM1[5018]<=26'd1993910; ROM2[5018]<=26'd11214468; ROM3[5018]<=26'd9750693; ROM4[5018]<=26'd23464727;
ROM1[5019]<=26'd1989809; ROM2[5019]<=26'd11213641; ROM3[5019]<=26'd9755446; ROM4[5019]<=26'd23464955;
ROM1[5020]<=26'd1991014; ROM2[5020]<=26'd11217798; ROM3[5020]<=26'd9764584; ROM4[5020]<=26'd23472507;
ROM1[5021]<=26'd1990291; ROM2[5021]<=26'd11220269; ROM3[5021]<=26'd9767694; ROM4[5021]<=26'd23475270;
ROM1[5022]<=26'd1991161; ROM2[5022]<=26'd11218437; ROM3[5022]<=26'd9760977; ROM4[5022]<=26'd23470441;
ROM1[5023]<=26'd2000379; ROM2[5023]<=26'd11218717; ROM3[5023]<=26'd9753237; ROM4[5023]<=26'd23468232;
ROM1[5024]<=26'd2002069; ROM2[5024]<=26'd11210825; ROM3[5024]<=26'd9739584; ROM4[5024]<=26'd23459380;
ROM1[5025]<=26'd1996451; ROM2[5025]<=26'd11208165; ROM3[5025]<=26'd9735650; ROM4[5025]<=26'd23455870;
ROM1[5026]<=26'd1991225; ROM2[5026]<=26'd11209412; ROM3[5026]<=26'd9739750; ROM4[5026]<=26'd23459345;
ROM1[5027]<=26'd1982531; ROM2[5027]<=26'd11205429; ROM3[5027]<=26'd9741351; ROM4[5027]<=26'd23458566;
ROM1[5028]<=26'd1975614; ROM2[5028]<=26'd11204079; ROM3[5028]<=26'd9743157; ROM4[5028]<=26'd23458077;
ROM1[5029]<=26'd1969894; ROM2[5029]<=26'd11199627; ROM3[5029]<=26'd9744100; ROM4[5029]<=26'd23455685;
ROM1[5030]<=26'd1973408; ROM2[5030]<=26'd11200932; ROM3[5030]<=26'd9742040; ROM4[5030]<=26'd23455135;
ROM1[5031]<=26'd1985735; ROM2[5031]<=26'd11205603; ROM3[5031]<=26'd9737873; ROM4[5031]<=26'd23456016;
ROM1[5032]<=26'd1999089; ROM2[5032]<=26'd11210397; ROM3[5032]<=26'd9735664; ROM4[5032]<=26'd23457320;
ROM1[5033]<=26'd2001336; ROM2[5033]<=26'd11213885; ROM3[5033]<=26'd9738559; ROM4[5033]<=26'd23462350;
ROM1[5034]<=26'd1993432; ROM2[5034]<=26'd11212230; ROM3[5034]<=26'd9741889; ROM4[5034]<=26'd23463362;
ROM1[5035]<=26'd1985680; ROM2[5035]<=26'd11210539; ROM3[5035]<=26'd9745875; ROM4[5035]<=26'd23462670;
ROM1[5036]<=26'd1981639; ROM2[5036]<=26'd11210804; ROM3[5036]<=26'd9749234; ROM4[5036]<=26'd23463807;
ROM1[5037]<=26'd1965804; ROM2[5037]<=26'd11200128; ROM3[5037]<=26'd9740373; ROM4[5037]<=26'd23452558;
ROM1[5038]<=26'd1961025; ROM2[5038]<=26'd11194662; ROM3[5038]<=26'd9736795; ROM4[5038]<=26'd23448621;
ROM1[5039]<=26'd1970033; ROM2[5039]<=26'd11199548; ROM3[5039]<=26'd9735765; ROM4[5039]<=26'd23451737;
ROM1[5040]<=26'd1980380; ROM2[5040]<=26'd11199614; ROM3[5040]<=26'd9727114; ROM4[5040]<=26'd23449822;
ROM1[5041]<=26'd1988025; ROM2[5041]<=26'd11202435; ROM3[5041]<=26'd9726559; ROM4[5041]<=26'd23451771;
ROM1[5042]<=26'd1985693; ROM2[5042]<=26'd11205727; ROM3[5042]<=26'd9730724; ROM4[5042]<=26'd23453290;
ROM1[5043]<=26'd1978723; ROM2[5043]<=26'd11203963; ROM3[5043]<=26'd9735347; ROM4[5043]<=26'd23454475;
ROM1[5044]<=26'd1972915; ROM2[5044]<=26'd11202417; ROM3[5044]<=26'd9738301; ROM4[5044]<=26'd23454539;
ROM1[5045]<=26'd1968977; ROM2[5045]<=26'd11203197; ROM3[5045]<=26'd9742169; ROM4[5045]<=26'd23456133;
ROM1[5046]<=26'd1969036; ROM2[5046]<=26'd11205439; ROM3[5046]<=26'd9746021; ROM4[5046]<=26'd23458618;
ROM1[5047]<=26'd1977295; ROM2[5047]<=26'd11210395; ROM3[5047]<=26'd9748173; ROM4[5047]<=26'd23463067;
ROM1[5048]<=26'd1992103; ROM2[5048]<=26'd11213937; ROM3[5048]<=26'd9746546; ROM4[5048]<=26'd23465072;
ROM1[5049]<=26'd1998662; ROM2[5049]<=26'd11210499; ROM3[5049]<=26'd9737757; ROM4[5049]<=26'd23461038;
ROM1[5050]<=26'd1992403; ROM2[5050]<=26'd11207116; ROM3[5050]<=26'd9733083; ROM4[5050]<=26'd23457088;
ROM1[5051]<=26'd1985791; ROM2[5051]<=26'd11208293; ROM3[5051]<=26'd9736082; ROM4[5051]<=26'd23458784;
ROM1[5052]<=26'd1973676; ROM2[5052]<=26'd11204759; ROM3[5052]<=26'd9734605; ROM4[5052]<=26'd23455584;
ROM1[5053]<=26'd1970494; ROM2[5053]<=26'd11205706; ROM3[5053]<=26'd9738897; ROM4[5053]<=26'd23457092;
ROM1[5054]<=26'd1973478; ROM2[5054]<=26'd11211102; ROM3[5054]<=26'd9748049; ROM4[5054]<=26'd23464799;
ROM1[5055]<=26'd1974576; ROM2[5055]<=26'd11210899; ROM3[5055]<=26'd9746815; ROM4[5055]<=26'd23463120;
ROM1[5056]<=26'd1979363; ROM2[5056]<=26'd11204189; ROM3[5056]<=26'd9737132; ROM4[5056]<=26'd23454115;
ROM1[5057]<=26'd1988193; ROM2[5057]<=26'd11202991; ROM3[5057]<=26'd9729780; ROM4[5057]<=26'd23453029;
ROM1[5058]<=26'd1989708; ROM2[5058]<=26'd11202737; ROM3[5058]<=26'd9729534; ROM4[5058]<=26'd23454048;
ROM1[5059]<=26'd1984592; ROM2[5059]<=26'd11200791; ROM3[5059]<=26'd9731811; ROM4[5059]<=26'd23452224;
ROM1[5060]<=26'd1981122; ROM2[5060]<=26'd11203083; ROM3[5060]<=26'd9739461; ROM4[5060]<=26'd23458373;
ROM1[5061]<=26'd1982164; ROM2[5061]<=26'd11207161; ROM3[5061]<=26'd9748874; ROM4[5061]<=26'd23464386;
ROM1[5062]<=26'd1975934; ROM2[5062]<=26'd11207469; ROM3[5062]<=26'd9752854; ROM4[5062]<=26'd23464767;
ROM1[5063]<=26'd1969332; ROM2[5063]<=26'd11201696; ROM3[5063]<=26'd9750403; ROM4[5063]<=26'd23461287;
ROM1[5064]<=26'd1978102; ROM2[5064]<=26'd11204559; ROM3[5064]<=26'd9749119; ROM4[5064]<=26'd23461469;
ROM1[5065]<=26'd1993360; ROM2[5065]<=26'd11210737; ROM3[5065]<=26'd9744178; ROM4[5065]<=26'd23463635;
ROM1[5066]<=26'd1999876; ROM2[5066]<=26'd11210550; ROM3[5066]<=26'd9741544; ROM4[5066]<=26'd23464114;
ROM1[5067]<=26'd1998425; ROM2[5067]<=26'd11212218; ROM3[5067]<=26'd9747123; ROM4[5067]<=26'd23466661;
ROM1[5068]<=26'd1990982; ROM2[5068]<=26'd11212295; ROM3[5068]<=26'd9751678; ROM4[5068]<=26'd23470085;
ROM1[5069]<=26'd1981773; ROM2[5069]<=26'd11207618; ROM3[5069]<=26'd9751016; ROM4[5069]<=26'd23466046;
ROM1[5070]<=26'd1975410; ROM2[5070]<=26'd11205685; ROM3[5070]<=26'd9751194; ROM4[5070]<=26'd23463674;
ROM1[5071]<=26'd1972420; ROM2[5071]<=26'd11205217; ROM3[5071]<=26'd9749638; ROM4[5071]<=26'd23462059;
ROM1[5072]<=26'd1976781; ROM2[5072]<=26'd11205717; ROM3[5072]<=26'd9746298; ROM4[5072]<=26'd23459744;
ROM1[5073]<=26'd1989998; ROM2[5073]<=26'd11208327; ROM3[5073]<=26'd9742677; ROM4[5073]<=26'd23460603;
ROM1[5074]<=26'd1997094; ROM2[5074]<=26'd11205279; ROM3[5074]<=26'd9732789; ROM4[5074]<=26'd23455747;
ROM1[5075]<=26'd1991050; ROM2[5075]<=26'd11201086; ROM3[5075]<=26'd9728050; ROM4[5075]<=26'd23451949;
ROM1[5076]<=26'd1986814; ROM2[5076]<=26'd11202426; ROM3[5076]<=26'd9733137; ROM4[5076]<=26'd23454609;
ROM1[5077]<=26'd1985293; ROM2[5077]<=26'd11205838; ROM3[5077]<=26'd9740653; ROM4[5077]<=26'd23458153;
ROM1[5078]<=26'd1977985; ROM2[5078]<=26'd11205499; ROM3[5078]<=26'd9742542; ROM4[5078]<=26'd23457973;
ROM1[5079]<=26'd1971047; ROM2[5079]<=26'd11202309; ROM3[5079]<=26'd9743308; ROM4[5079]<=26'd23457582;
ROM1[5080]<=26'd1972996; ROM2[5080]<=26'd11202584; ROM3[5080]<=26'd9742354; ROM4[5080]<=26'd23457341;
ROM1[5081]<=26'd1980638; ROM2[5081]<=26'd11203909; ROM3[5081]<=26'd9738055; ROM4[5081]<=26'd23456507;
ROM1[5082]<=26'd1993097; ROM2[5082]<=26'd11202934; ROM3[5082]<=26'd9733012; ROM4[5082]<=26'd23454242;
ROM1[5083]<=26'd1995834; ROM2[5083]<=26'd11204689; ROM3[5083]<=26'd9732807; ROM4[5083]<=26'd23454515;
ROM1[5084]<=26'd1991115; ROM2[5084]<=26'd11207747; ROM3[5084]<=26'd9736053; ROM4[5084]<=26'd23457171;
ROM1[5085]<=26'd1985912; ROM2[5085]<=26'd11208192; ROM3[5085]<=26'd9738580; ROM4[5085]<=26'd23458109;
ROM1[5086]<=26'd1981891; ROM2[5086]<=26'd11210803; ROM3[5086]<=26'd9742846; ROM4[5086]<=26'd23462212;
ROM1[5087]<=26'd1969120; ROM2[5087]<=26'd11202328; ROM3[5087]<=26'd9739810; ROM4[5087]<=26'd23455321;
ROM1[5088]<=26'd1960090; ROM2[5088]<=26'd11193002; ROM3[5088]<=26'd9735370; ROM4[5088]<=26'd23446893;
ROM1[5089]<=26'd1967725; ROM2[5089]<=26'd11195022; ROM3[5089]<=26'd9736154; ROM4[5089]<=26'd23448853;
ROM1[5090]<=26'd1979256; ROM2[5090]<=26'd11194157; ROM3[5090]<=26'd9729885; ROM4[5090]<=26'd23447174;
ROM1[5091]<=26'd1986280; ROM2[5091]<=26'd11195852; ROM3[5091]<=26'd9726993; ROM4[5091]<=26'd23448579;
ROM1[5092]<=26'd1986725; ROM2[5092]<=26'd11199462; ROM3[5092]<=26'd9731460; ROM4[5092]<=26'd23452517;
ROM1[5093]<=26'd1975370; ROM2[5093]<=26'd11193816; ROM3[5093]<=26'd9731224; ROM4[5093]<=26'd23448106;
ROM1[5094]<=26'd1965198; ROM2[5094]<=26'd11189538; ROM3[5094]<=26'd9732110; ROM4[5094]<=26'd23445635;
ROM1[5095]<=26'd1960912; ROM2[5095]<=26'd11189228; ROM3[5095]<=26'd9737394; ROM4[5095]<=26'd23448107;
ROM1[5096]<=26'd1957664; ROM2[5096]<=26'd11187696; ROM3[5096]<=26'd9739457; ROM4[5096]<=26'd23449320;
ROM1[5097]<=26'd1963786; ROM2[5097]<=26'd11188415; ROM3[5097]<=26'd9740346; ROM4[5097]<=26'd23452325;
ROM1[5098]<=26'd1981009; ROM2[5098]<=26'd11194941; ROM3[5098]<=26'd9741461; ROM4[5098]<=26'd23457047;
ROM1[5099]<=26'd1993874; ROM2[5099]<=26'd11201791; ROM3[5099]<=26'd9740632; ROM4[5099]<=26'd23460456;
ROM1[5100]<=26'd1992778; ROM2[5100]<=26'd11202993; ROM3[5100]<=26'd9739533; ROM4[5100]<=26'd23460485;
ROM1[5101]<=26'd1989593; ROM2[5101]<=26'd11207133; ROM3[5101]<=26'd9744732; ROM4[5101]<=26'd23464067;
ROM1[5102]<=26'd1988638; ROM2[5102]<=26'd11209785; ROM3[5102]<=26'd9751584; ROM4[5102]<=26'd23467549;
ROM1[5103]<=26'd1977292; ROM2[5103]<=26'd11202134; ROM3[5103]<=26'd9746951; ROM4[5103]<=26'd23460725;
ROM1[5104]<=26'd1968397; ROM2[5104]<=26'd11197818; ROM3[5104]<=26'd9743636; ROM4[5104]<=26'd23455565;
ROM1[5105]<=26'd1972780; ROM2[5105]<=26'd11199336; ROM3[5105]<=26'd9742449; ROM4[5105]<=26'd23456662;
ROM1[5106]<=26'd1982913; ROM2[5106]<=26'd11200676; ROM3[5106]<=26'd9737688; ROM4[5106]<=26'd23457169;
ROM1[5107]<=26'd2000964; ROM2[5107]<=26'd11206377; ROM3[5107]<=26'd9737456; ROM4[5107]<=26'd23462692;
ROM1[5108]<=26'd1999351; ROM2[5108]<=26'd11201824; ROM3[5108]<=26'd9736113; ROM4[5108]<=26'd23459448;
ROM1[5109]<=26'd1982542; ROM2[5109]<=26'd11190705; ROM3[5109]<=26'd9731998; ROM4[5109]<=26'd23450676;
ROM1[5110]<=26'd1972451; ROM2[5110]<=26'd11187544; ROM3[5110]<=26'd9734618; ROM4[5110]<=26'd23449691;
ROM1[5111]<=26'd1969257; ROM2[5111]<=26'd11188068; ROM3[5111]<=26'd9738704; ROM4[5111]<=26'd23451144;
ROM1[5112]<=26'd1964932; ROM2[5112]<=26'd11190209; ROM3[5112]<=26'd9742345; ROM4[5112]<=26'd23453760;
ROM1[5113]<=26'd1968246; ROM2[5113]<=26'd11193428; ROM3[5113]<=26'd9748153; ROM4[5113]<=26'd23457342;
ROM1[5114]<=26'd1975939; ROM2[5114]<=26'd11195533; ROM3[5114]<=26'd9747487; ROM4[5114]<=26'd23459394;
ROM1[5115]<=26'd1985429; ROM2[5115]<=26'd11194659; ROM3[5115]<=26'd9739635; ROM4[5115]<=26'd23458541;
ROM1[5116]<=26'd1989781; ROM2[5116]<=26'd11191915; ROM3[5116]<=26'd9735289; ROM4[5116]<=26'd23456555;
ROM1[5117]<=26'd1986150; ROM2[5117]<=26'd11192846; ROM3[5117]<=26'd9738360; ROM4[5117]<=26'd23457923;
ROM1[5118]<=26'd1980854; ROM2[5118]<=26'd11195018; ROM3[5118]<=26'd9745514; ROM4[5118]<=26'd23461507;
ROM1[5119]<=26'd1976777; ROM2[5119]<=26'd11196430; ROM3[5119]<=26'd9751523; ROM4[5119]<=26'd23462774;
ROM1[5120]<=26'd1972060; ROM2[5120]<=26'd11196770; ROM3[5120]<=26'd9752688; ROM4[5120]<=26'd23463802;
ROM1[5121]<=26'd1966687; ROM2[5121]<=26'd11195993; ROM3[5121]<=26'd9747878; ROM4[5121]<=26'd23460792;
ROM1[5122]<=26'd1967842; ROM2[5122]<=26'd11193414; ROM3[5122]<=26'd9741227; ROM4[5122]<=26'd23454705;
ROM1[5123]<=26'd1980860; ROM2[5123]<=26'd11194477; ROM3[5123]<=26'd9737028; ROM4[5123]<=26'd23454722;
ROM1[5124]<=26'd1991320; ROM2[5124]<=26'd11195529; ROM3[5124]<=26'd9735155; ROM4[5124]<=26'd23455366;
ROM1[5125]<=26'd1988285; ROM2[5125]<=26'd11193024; ROM3[5125]<=26'd9738027; ROM4[5125]<=26'd23455754;
ROM1[5126]<=26'd1979087; ROM2[5126]<=26'd11191131; ROM3[5126]<=26'd9738493; ROM4[5126]<=26'd23454178;
ROM1[5127]<=26'd1972597; ROM2[5127]<=26'd11191364; ROM3[5127]<=26'd9742745; ROM4[5127]<=26'd23455022;
ROM1[5128]<=26'd1970038; ROM2[5128]<=26'd11192715; ROM3[5128]<=26'd9749285; ROM4[5128]<=26'd23460770;
ROM1[5129]<=26'd1969797; ROM2[5129]<=26'd11196521; ROM3[5129]<=26'd9755913; ROM4[5129]<=26'd23465361;
ROM1[5130]<=26'd1972688; ROM2[5130]<=26'd11197620; ROM3[5130]<=26'd9757968; ROM4[5130]<=26'd23467968;
ROM1[5131]<=26'd1979723; ROM2[5131]<=26'd11195501; ROM3[5131]<=26'd9750677; ROM4[5131]<=26'd23464762;
ROM1[5132]<=26'd1992173; ROM2[5132]<=26'd11196175; ROM3[5132]<=26'd9744632; ROM4[5132]<=26'd23462489;
ROM1[5133]<=26'd1994945; ROM2[5133]<=26'd11196350; ROM3[5133]<=26'd9743204; ROM4[5133]<=26'd23463231;
ROM1[5134]<=26'd1989581; ROM2[5134]<=26'd11197107; ROM3[5134]<=26'd9745598; ROM4[5134]<=26'd23464396;
ROM1[5135]<=26'd1981203; ROM2[5135]<=26'd11196690; ROM3[5135]<=26'd9747701; ROM4[5135]<=26'd23462803;
ROM1[5136]<=26'd1979081; ROM2[5136]<=26'd11199436; ROM3[5136]<=26'd9752446; ROM4[5136]<=26'd23465288;
ROM1[5137]<=26'd1973419; ROM2[5137]<=26'd11200861; ROM3[5137]<=26'd9754205; ROM4[5137]<=26'd23465752;
ROM1[5138]<=26'd1971638; ROM2[5138]<=26'd11199144; ROM3[5138]<=26'd9751159; ROM4[5138]<=26'd23463073;
ROM1[5139]<=26'd1981988; ROM2[5139]<=26'd11202893; ROM3[5139]<=26'd9752861; ROM4[5139]<=26'd23465526;
ROM1[5140]<=26'd2003752; ROM2[5140]<=26'd11214528; ROM3[5140]<=26'd9756332; ROM4[5140]<=26'd23474146;
ROM1[5141]<=26'd2013415; ROM2[5141]<=26'd11218925; ROM3[5141]<=26'd9756108; ROM4[5141]<=26'd23477235;
ROM1[5142]<=26'd1993791; ROM2[5142]<=26'd11203911; ROM3[5142]<=26'd9744243; ROM4[5142]<=26'd23461677;
ROM1[5143]<=26'd1982134; ROM2[5143]<=26'd11199200; ROM3[5143]<=26'd9740764; ROM4[5143]<=26'd23456818;
ROM1[5144]<=26'd1975786; ROM2[5144]<=26'd11199622; ROM3[5144]<=26'd9742839; ROM4[5144]<=26'd23456045;
ROM1[5145]<=26'd1968991; ROM2[5145]<=26'd11197019; ROM3[5145]<=26'd9742372; ROM4[5145]<=26'd23453607;
ROM1[5146]<=26'd1975767; ROM2[5146]<=26'd11204692; ROM3[5146]<=26'd9751073; ROM4[5146]<=26'd23462521;
ROM1[5147]<=26'd1981780; ROM2[5147]<=26'd11207487; ROM3[5147]<=26'd9751062; ROM4[5147]<=26'd23464517;
ROM1[5148]<=26'd1986465; ROM2[5148]<=26'd11203303; ROM3[5148]<=26'd9737649; ROM4[5148]<=26'd23455890;
ROM1[5149]<=26'd1995193; ROM2[5149]<=26'd11203733; ROM3[5149]<=26'd9732753; ROM4[5149]<=26'd23455483;
ROM1[5150]<=26'd1994776; ROM2[5150]<=26'd11204344; ROM3[5150]<=26'd9735787; ROM4[5150]<=26'd23457829;
ROM1[5151]<=26'd1984293; ROM2[5151]<=26'd11199679; ROM3[5151]<=26'd9735944; ROM4[5151]<=26'd23454574;
ROM1[5152]<=26'd1981454; ROM2[5152]<=26'd11204083; ROM3[5152]<=26'd9745080; ROM4[5152]<=26'd23460812;
ROM1[5153]<=26'd1969421; ROM2[5153]<=26'd11199580; ROM3[5153]<=26'd9742641; ROM4[5153]<=26'd23456590;
ROM1[5154]<=26'd1951156; ROM2[5154]<=26'd11187434; ROM3[5154]<=26'd9729674; ROM4[5154]<=26'd23444171;
ROM1[5155]<=26'd1951809; ROM2[5155]<=26'd11186727; ROM3[5155]<=26'd9726914; ROM4[5155]<=26'd23442661;
ROM1[5156]<=26'd1959517; ROM2[5156]<=26'd11183378; ROM3[5156]<=26'd9720077; ROM4[5156]<=26'd23439424;
ROM1[5157]<=26'd1976715; ROM2[5157]<=26'd11184343; ROM3[5157]<=26'd9715620; ROM4[5157]<=26'd23438784;
ROM1[5158]<=26'd1989503; ROM2[5158]<=26'd11193047; ROM3[5158]<=26'd9725568; ROM4[5158]<=26'd23448267;
ROM1[5159]<=26'd1986476; ROM2[5159]<=26'd11194311; ROM3[5159]<=26'd9733558; ROM4[5159]<=26'd23454124;
ROM1[5160]<=26'd1973888; ROM2[5160]<=26'd11186612; ROM3[5160]<=26'd9735184; ROM4[5160]<=26'd23452210;
ROM1[5161]<=26'd1965793; ROM2[5161]<=26'd11184035; ROM3[5161]<=26'd9737275; ROM4[5161]<=26'd23450589;
ROM1[5162]<=26'd1961254; ROM2[5162]<=26'd11184684; ROM3[5162]<=26'd9740381; ROM4[5162]<=26'd23450883;
ROM1[5163]<=26'd1961649; ROM2[5163]<=26'd11184905; ROM3[5163]<=26'd9739913; ROM4[5163]<=26'd23451317;
ROM1[5164]<=26'd1970203; ROM2[5164]<=26'd11186286; ROM3[5164]<=26'd9737583; ROM4[5164]<=26'd23451088;
ROM1[5165]<=26'd1982195; ROM2[5165]<=26'd11187244; ROM3[5165]<=26'd9734020; ROM4[5165]<=26'd23452126;
ROM1[5166]<=26'd1987882; ROM2[5166]<=26'd11188709; ROM3[5166]<=26'd9735329; ROM4[5166]<=26'd23454138;
ROM1[5167]<=26'd1985764; ROM2[5167]<=26'd11189678; ROM3[5167]<=26'd9738902; ROM4[5167]<=26'd23455843;
ROM1[5168]<=26'd1980674; ROM2[5168]<=26'd11189881; ROM3[5168]<=26'd9741323; ROM4[5168]<=26'd23455189;
ROM1[5169]<=26'd1978395; ROM2[5169]<=26'd11191565; ROM3[5169]<=26'd9745673; ROM4[5169]<=26'd23457085;
ROM1[5170]<=26'd1975804; ROM2[5170]<=26'd11193547; ROM3[5170]<=26'd9747836; ROM4[5170]<=26'd23459231;
ROM1[5171]<=26'd1970909; ROM2[5171]<=26'd11192422; ROM3[5171]<=26'd9749117; ROM4[5171]<=26'd23457776;
ROM1[5172]<=26'd1980601; ROM2[5172]<=26'd11198086; ROM3[5172]<=26'd9753861; ROM4[5172]<=26'd23463434;
ROM1[5173]<=26'd1993024; ROM2[5173]<=26'd11199955; ROM3[5173]<=26'd9751424; ROM4[5173]<=26'd23464582;
ROM1[5174]<=26'd1999436; ROM2[5174]<=26'd11196669; ROM3[5174]<=26'd9745043; ROM4[5174]<=26'd23460544;
ROM1[5175]<=26'd2001416; ROM2[5175]<=26'd11198052; ROM3[5175]<=26'd9747700; ROM4[5175]<=26'd23462443;
ROM1[5176]<=26'd1991850; ROM2[5176]<=26'd11194754; ROM3[5176]<=26'd9748497; ROM4[5176]<=26'd23461435;
ROM1[5177]<=26'd1981558; ROM2[5177]<=26'd11188733; ROM3[5177]<=26'd9747952; ROM4[5177]<=26'd23457537;
ROM1[5178]<=26'd1976775; ROM2[5178]<=26'd11190089; ROM3[5178]<=26'd9751475; ROM4[5178]<=26'd23461112;
ROM1[5179]<=26'd1971830; ROM2[5179]<=26'd11190448; ROM3[5179]<=26'd9752950; ROM4[5179]<=26'd23463003;
ROM1[5180]<=26'd1973614; ROM2[5180]<=26'd11190042; ROM3[5180]<=26'd9752042; ROM4[5180]<=26'd23462333;
ROM1[5181]<=26'd1987753; ROM2[5181]<=26'd11196105; ROM3[5181]<=26'd9750961; ROM4[5181]<=26'd23467877;
ROM1[5182]<=26'd2002676; ROM2[5182]<=26'd11198799; ROM3[5182]<=26'd9748527; ROM4[5182]<=26'd23469096;
ROM1[5183]<=26'd2002112; ROM2[5183]<=26'd11198421; ROM3[5183]<=26'd9747583; ROM4[5183]<=26'd23468307;
ROM1[5184]<=26'd1995363; ROM2[5184]<=26'd11197315; ROM3[5184]<=26'd9748979; ROM4[5184]<=26'd23467811;
ROM1[5185]<=26'd1993539; ROM2[5185]<=26'd11200653; ROM3[5185]<=26'd9755137; ROM4[5185]<=26'd23470805;
ROM1[5186]<=26'd1993839; ROM2[5186]<=26'd11204454; ROM3[5186]<=26'd9762814; ROM4[5186]<=26'd23475000;
ROM1[5187]<=26'd1987145; ROM2[5187]<=26'd11202956; ROM3[5187]<=26'd9766149; ROM4[5187]<=26'd23474581;
ROM1[5188]<=26'd1979765; ROM2[5188]<=26'd11195809; ROM3[5188]<=26'd9759729; ROM4[5188]<=26'd23467982;
ROM1[5189]<=26'd1976800; ROM2[5189]<=26'd11187152; ROM3[5189]<=26'd9747398; ROM4[5189]<=26'd23458079;
ROM1[5190]<=26'd1985229; ROM2[5190]<=26'd11184254; ROM3[5190]<=26'd9737082; ROM4[5190]<=26'd23451992;
ROM1[5191]<=26'd1992873; ROM2[5191]<=26'd11186643; ROM3[5191]<=26'd9733350; ROM4[5191]<=26'd23452066;
ROM1[5192]<=26'd1993371; ROM2[5192]<=26'd11192201; ROM3[5192]<=26'd9738693; ROM4[5192]<=26'd23456458;
ROM1[5193]<=26'd1989494; ROM2[5193]<=26'd11195052; ROM3[5193]<=26'd9747745; ROM4[5193]<=26'd23460753;
ROM1[5194]<=26'd1982948; ROM2[5194]<=26'd11193761; ROM3[5194]<=26'd9750766; ROM4[5194]<=26'd23461710;
ROM1[5195]<=26'd1973886; ROM2[5195]<=26'd11190206; ROM3[5195]<=26'd9748785; ROM4[5195]<=26'd23457614;
ROM1[5196]<=26'd1970924; ROM2[5196]<=26'd11191603; ROM3[5196]<=26'd9748484; ROM4[5196]<=26'd23457597;
ROM1[5197]<=26'd1977809; ROM2[5197]<=26'd11193796; ROM3[5197]<=26'd9748340; ROM4[5197]<=26'd23458746;
ROM1[5198]<=26'd1994610; ROM2[5198]<=26'd11200079; ROM3[5198]<=26'd9748584; ROM4[5198]<=26'd23463775;
ROM1[5199]<=26'd2010172; ROM2[5199]<=26'd11204812; ROM3[5199]<=26'd9747780; ROM4[5199]<=26'd23467930;
ROM1[5200]<=26'd1992823; ROM2[5200]<=26'd11189570; ROM3[5200]<=26'd9732657; ROM4[5200]<=26'd23453023;
ROM1[5201]<=26'd1975543; ROM2[5201]<=26'd11181695; ROM3[5201]<=26'd9726696; ROM4[5201]<=26'd23446763;
ROM1[5202]<=26'd1968941; ROM2[5202]<=26'd11179606; ROM3[5202]<=26'd9728800; ROM4[5202]<=26'd23446370;
ROM1[5203]<=26'd1961295; ROM2[5203]<=26'd11177279; ROM3[5203]<=26'd9730093; ROM4[5203]<=26'd23446624;
ROM1[5204]<=26'd1965366; ROM2[5204]<=26'd11183445; ROM3[5204]<=26'd9739645; ROM4[5204]<=26'd23455573;
ROM1[5205]<=26'd1965736; ROM2[5205]<=26'd11180481; ROM3[5205]<=26'd9735666; ROM4[5205]<=26'd23450634;
ROM1[5206]<=26'd1965876; ROM2[5206]<=26'd11174051; ROM3[5206]<=26'd9724184; ROM4[5206]<=26'd23441027;
ROM1[5207]<=26'd1978875; ROM2[5207]<=26'd11174738; ROM3[5207]<=26'd9721434; ROM4[5207]<=26'd23442506;
ROM1[5208]<=26'd1985875; ROM2[5208]<=26'd11176973; ROM3[5208]<=26'd9727480; ROM4[5208]<=26'd23449090;
ROM1[5209]<=26'd1981813; ROM2[5209]<=26'd11181394; ROM3[5209]<=26'd9735469; ROM4[5209]<=26'd23453894;
ROM1[5210]<=26'd1975219; ROM2[5210]<=26'd11183086; ROM3[5210]<=26'd9739552; ROM4[5210]<=26'd23455965;
ROM1[5211]<=26'd1972881; ROM2[5211]<=26'd11185120; ROM3[5211]<=26'd9742695; ROM4[5211]<=26'd23458333;
ROM1[5212]<=26'd1970866; ROM2[5212]<=26'd11189712; ROM3[5212]<=26'd9748320; ROM4[5212]<=26'd23461413;
ROM1[5213]<=26'd1968513; ROM2[5213]<=26'd11184379; ROM3[5213]<=26'd9746344; ROM4[5213]<=26'd23458809;
ROM1[5214]<=26'd1976301; ROM2[5214]<=26'd11184395; ROM3[5214]<=26'd9744486; ROM4[5214]<=26'd23458990;
ROM1[5215]<=26'd1985632; ROM2[5215]<=26'd11185748; ROM3[5215]<=26'd9737096; ROM4[5215]<=26'd23455870;
ROM1[5216]<=26'd1984424; ROM2[5216]<=26'd11181410; ROM3[5216]<=26'd9727280; ROM4[5216]<=26'd23448526;
ROM1[5217]<=26'd1982429; ROM2[5217]<=26'd11182617; ROM3[5217]<=26'd9729383; ROM4[5217]<=26'd23451056;
ROM1[5218]<=26'd1976126; ROM2[5218]<=26'd11180820; ROM3[5218]<=26'd9734111; ROM4[5218]<=26'd23452890;
ROM1[5219]<=26'd1968530; ROM2[5219]<=26'd11178005; ROM3[5219]<=26'd9736581; ROM4[5219]<=26'd23452661;
ROM1[5220]<=26'd1962400; ROM2[5220]<=26'd11178675; ROM3[5220]<=26'd9741531; ROM4[5220]<=26'd23455321;
ROM1[5221]<=26'd1960761; ROM2[5221]<=26'd11180555; ROM3[5221]<=26'd9745471; ROM4[5221]<=26'd23456214;
ROM1[5222]<=26'd1967012; ROM2[5222]<=26'd11181468; ROM3[5222]<=26'd9745246; ROM4[5222]<=26'd23456570;
ROM1[5223]<=26'd1979822; ROM2[5223]<=26'd11181094; ROM3[5223]<=26'd9741429; ROM4[5223]<=26'd23456384;
ROM1[5224]<=26'd1992798; ROM2[5224]<=26'd11182988; ROM3[5224]<=26'd9741337; ROM4[5224]<=26'd23459857;
ROM1[5225]<=26'd1992457; ROM2[5225]<=26'd11184828; ROM3[5225]<=26'd9743273; ROM4[5225]<=26'd23462624;
ROM1[5226]<=26'd1986610; ROM2[5226]<=26'd11186097; ROM3[5226]<=26'd9747763; ROM4[5226]<=26'd23464808;
ROM1[5227]<=26'd1977824; ROM2[5227]<=26'd11183252; ROM3[5227]<=26'd9749508; ROM4[5227]<=26'd23462759;
ROM1[5228]<=26'd1972279; ROM2[5228]<=26'd11182413; ROM3[5228]<=26'd9750702; ROM4[5228]<=26'd23462625;
ROM1[5229]<=26'd1970488; ROM2[5229]<=26'd11182604; ROM3[5229]<=26'd9755733; ROM4[5229]<=26'd23466322;
ROM1[5230]<=26'd1973379; ROM2[5230]<=26'd11183387; ROM3[5230]<=26'd9755573; ROM4[5230]<=26'd23468157;
ROM1[5231]<=26'd1984081; ROM2[5231]<=26'd11183578; ROM3[5231]<=26'd9754744; ROM4[5231]<=26'd23468509;
ROM1[5232]<=26'd1990998; ROM2[5232]<=26'd11179294; ROM3[5232]<=26'd9747043; ROM4[5232]<=26'd23462803;
ROM1[5233]<=26'd1989652; ROM2[5233]<=26'd11178303; ROM3[5233]<=26'd9744785; ROM4[5233]<=26'd23461668;
ROM1[5234]<=26'd1978024; ROM2[5234]<=26'd11172962; ROM3[5234]<=26'd9743025; ROM4[5234]<=26'd23458225;
ROM1[5235]<=26'd1966215; ROM2[5235]<=26'd11168478; ROM3[5235]<=26'd9740042; ROM4[5235]<=26'd23454186;
ROM1[5236]<=26'd1965182; ROM2[5236]<=26'd11170453; ROM3[5236]<=26'd9742684; ROM4[5236]<=26'd23455512;
ROM1[5237]<=26'd1959030; ROM2[5237]<=26'd11168895; ROM3[5237]<=26'd9742597; ROM4[5237]<=26'd23453236;
ROM1[5238]<=26'd1955566; ROM2[5238]<=26'd11166789; ROM3[5238]<=26'd9739839; ROM4[5238]<=26'd23450943;
ROM1[5239]<=26'd1966812; ROM2[5239]<=26'd11170970; ROM3[5239]<=26'd9742216; ROM4[5239]<=26'd23456897;
ROM1[5240]<=26'd1981454; ROM2[5240]<=26'd11173247; ROM3[5240]<=26'd9741429; ROM4[5240]<=26'd23458984;
ROM1[5241]<=26'd1984845; ROM2[5241]<=26'd11172495; ROM3[5241]<=26'd9736083; ROM4[5241]<=26'd23455855;
ROM1[5242]<=26'd1979791; ROM2[5242]<=26'd11170924; ROM3[5242]<=26'd9734858; ROM4[5242]<=26'd23454213;
ROM1[5243]<=26'd1971201; ROM2[5243]<=26'd11168338; ROM3[5243]<=26'd9735681; ROM4[5243]<=26'd23450757;
ROM1[5244]<=26'd1959875; ROM2[5244]<=26'd11163335; ROM3[5244]<=26'd9735633; ROM4[5244]<=26'd23448210;
ROM1[5245]<=26'd1954441; ROM2[5245]<=26'd11161723; ROM3[5245]<=26'd9738257; ROM4[5245]<=26'd23450191;
ROM1[5246]<=26'd1954185; ROM2[5246]<=26'd11165508; ROM3[5246]<=26'd9741683; ROM4[5246]<=26'd23451795;
ROM1[5247]<=26'd1958029; ROM2[5247]<=26'd11166908; ROM3[5247]<=26'd9738254; ROM4[5247]<=26'd23450515;
ROM1[5248]<=26'd1970137; ROM2[5248]<=26'd11170737; ROM3[5248]<=26'd9732385; ROM4[5248]<=26'd23450656;
ROM1[5249]<=26'd1979768; ROM2[5249]<=26'd11174281; ROM3[5249]<=26'd9731555; ROM4[5249]<=26'd23452123;
ROM1[5250]<=26'd1980723; ROM2[5250]<=26'd11175970; ROM3[5250]<=26'd9735831; ROM4[5250]<=26'd23454336;
ROM1[5251]<=26'd1975406; ROM2[5251]<=26'd11177951; ROM3[5251]<=26'd9739411; ROM4[5251]<=26'd23455022;
ROM1[5252]<=26'd1977868; ROM2[5252]<=26'd11187374; ROM3[5252]<=26'd9750113; ROM4[5252]<=26'd23463513;
ROM1[5253]<=26'd1978826; ROM2[5253]<=26'd11192463; ROM3[5253]<=26'd9757541; ROM4[5253]<=26'd23469405;
ROM1[5254]<=26'd1962823; ROM2[5254]<=26'd11180211; ROM3[5254]<=26'd9748958; ROM4[5254]<=26'd23458311;
ROM1[5255]<=26'd1953897; ROM2[5255]<=26'd11169417; ROM3[5255]<=26'd9739543; ROM4[5255]<=26'd23448423;
ROM1[5256]<=26'd1958099; ROM2[5256]<=26'd11165066; ROM3[5256]<=26'd9730372; ROM4[5256]<=26'd23443266;
ROM1[5257]<=26'd1967219; ROM2[5257]<=26'd11163998; ROM3[5257]<=26'd9721278; ROM4[5257]<=26'd23439790;
ROM1[5258]<=26'd1972737; ROM2[5258]<=26'd11168676; ROM3[5258]<=26'd9722942; ROM4[5258]<=26'd23443883;
ROM1[5259]<=26'd1972788; ROM2[5259]<=26'd11175085; ROM3[5259]<=26'd9731718; ROM4[5259]<=26'd23449568;
ROM1[5260]<=26'd1963294; ROM2[5260]<=26'd11172398; ROM3[5260]<=26'd9733092; ROM4[5260]<=26'd23446080;
ROM1[5261]<=26'd1955127; ROM2[5261]<=26'd11167116; ROM3[5261]<=26'd9729410; ROM4[5261]<=26'd23441146;
ROM1[5262]<=26'd1952042; ROM2[5262]<=26'd11169031; ROM3[5262]<=26'd9732284; ROM4[5262]<=26'd23444160;
ROM1[5263]<=26'd1953415; ROM2[5263]<=26'd11170495; ROM3[5263]<=26'd9733888; ROM4[5263]<=26'd23445056;
ROM1[5264]<=26'd1959951; ROM2[5264]<=26'd11170051; ROM3[5264]<=26'd9730246; ROM4[5264]<=26'd23442711;
ROM1[5265]<=26'd1971416; ROM2[5265]<=26'd11171144; ROM3[5265]<=26'd9724346; ROM4[5265]<=26'd23440454;
ROM1[5266]<=26'd1976651; ROM2[5266]<=26'd11170628; ROM3[5266]<=26'd9722679; ROM4[5266]<=26'd23440859;
ROM1[5267]<=26'd1973364; ROM2[5267]<=26'd11170358; ROM3[5267]<=26'd9724912; ROM4[5267]<=26'd23443181;
ROM1[5268]<=26'd1969070; ROM2[5268]<=26'd11171308; ROM3[5268]<=26'd9729874; ROM4[5268]<=26'd23445551;
ROM1[5269]<=26'd1969978; ROM2[5269]<=26'd11175128; ROM3[5269]<=26'd9740644; ROM4[5269]<=26'd23451188;
ROM1[5270]<=26'd1966736; ROM2[5270]<=26'd11177597; ROM3[5270]<=26'd9747478; ROM4[5270]<=26'd23453141;
ROM1[5271]<=26'd1962324; ROM2[5271]<=26'd11176142; ROM3[5271]<=26'd9746151; ROM4[5271]<=26'd23451456;
ROM1[5272]<=26'd1956677; ROM2[5272]<=26'd11165271; ROM3[5272]<=26'd9734098; ROM4[5272]<=26'd23441206;
ROM1[5273]<=26'd1958760; ROM2[5273]<=26'd11156281; ROM3[5273]<=26'd9720352; ROM4[5273]<=26'd23431777;
ROM1[5274]<=26'd1969071; ROM2[5274]<=26'd11159713; ROM3[5274]<=26'd9716344; ROM4[5274]<=26'd23432036;
ROM1[5275]<=26'd1968225; ROM2[5275]<=26'd11161430; ROM3[5275]<=26'd9719709; ROM4[5275]<=26'd23434373;
ROM1[5276]<=26'd1967281; ROM2[5276]<=26'd11166200; ROM3[5276]<=26'd9725384; ROM4[5276]<=26'd23437636;
ROM1[5277]<=26'd1961895; ROM2[5277]<=26'd11167335; ROM3[5277]<=26'd9727948; ROM4[5277]<=26'd23437918;
ROM1[5278]<=26'd1954633; ROM2[5278]<=26'd11163922; ROM3[5278]<=26'd9727664; ROM4[5278]<=26'd23436253;
ROM1[5279]<=26'd1950318; ROM2[5279]<=26'd11163171; ROM3[5279]<=26'd9729855; ROM4[5279]<=26'd23435685;
ROM1[5280]<=26'd1951841; ROM2[5280]<=26'd11165092; ROM3[5280]<=26'd9732532; ROM4[5280]<=26'd23437515;
ROM1[5281]<=26'd1965852; ROM2[5281]<=26'd11169441; ROM3[5281]<=26'd9733495; ROM4[5281]<=26'd23441497;
ROM1[5282]<=26'd1980770; ROM2[5282]<=26'd11172885; ROM3[5282]<=26'd9730123; ROM4[5282]<=26'd23443822;
ROM1[5283]<=26'd1980408; ROM2[5283]<=26'd11170953; ROM3[5283]<=26'd9726806; ROM4[5283]<=26'd23441970;
ROM1[5284]<=26'd1974923; ROM2[5284]<=26'd11172744; ROM3[5284]<=26'd9731637; ROM4[5284]<=26'd23445094;
ROM1[5285]<=26'd1973973; ROM2[5285]<=26'd11179544; ROM3[5285]<=26'd9743103; ROM4[5285]<=26'd23452837;
ROM1[5286]<=26'd1967467; ROM2[5286]<=26'd11175907; ROM3[5286]<=26'd9742646; ROM4[5286]<=26'd23449439;
ROM1[5287]<=26'd1957516; ROM2[5287]<=26'd11170363; ROM3[5287]<=26'd9738178; ROM4[5287]<=26'd23443859;
ROM1[5288]<=26'd1958258; ROM2[5288]<=26'd11170281; ROM3[5288]<=26'd9737690; ROM4[5288]<=26'd23445007;
ROM1[5289]<=26'd1960870; ROM2[5289]<=26'd11166441; ROM3[5289]<=26'd9728906; ROM4[5289]<=26'd23441238;
ROM1[5290]<=26'd1970931; ROM2[5290]<=26'd11165818; ROM3[5290]<=26'd9723113; ROM4[5290]<=26'd23438841;
ROM1[5291]<=26'd1978692; ROM2[5291]<=26'd11169800; ROM3[5291]<=26'd9724088; ROM4[5291]<=26'd23442878;
ROM1[5292]<=26'd1976078; ROM2[5292]<=26'd11170345; ROM3[5292]<=26'd9728592; ROM4[5292]<=26'd23445044;
ROM1[5293]<=26'd1967103; ROM2[5293]<=26'd11167935; ROM3[5293]<=26'd9731625; ROM4[5293]<=26'd23444582;
ROM1[5294]<=26'd1964418; ROM2[5294]<=26'd11170869; ROM3[5294]<=26'd9738196; ROM4[5294]<=26'd23450060;
ROM1[5295]<=26'd1964998; ROM2[5295]<=26'd11176322; ROM3[5295]<=26'd9747062; ROM4[5295]<=26'd23457698;
ROM1[5296]<=26'd1960116; ROM2[5296]<=26'd11173337; ROM3[5296]<=26'd9744280; ROM4[5296]<=26'd23454787;
ROM1[5297]<=26'd1961553; ROM2[5297]<=26'd11168751; ROM3[5297]<=26'd9739197; ROM4[5297]<=26'd23450214;
ROM1[5298]<=26'd1976260; ROM2[5298]<=26'd11172187; ROM3[5298]<=26'd9736928; ROM4[5298]<=26'd23453115;
ROM1[5299]<=26'd1988402; ROM2[5299]<=26'd11174589; ROM3[5299]<=26'd9734605; ROM4[5299]<=26'd23454913;
ROM1[5300]<=26'd1987042; ROM2[5300]<=26'd11174439; ROM3[5300]<=26'd9736180; ROM4[5300]<=26'd23455494;
ROM1[5301]<=26'd1979822; ROM2[5301]<=26'd11174946; ROM3[5301]<=26'd9738700; ROM4[5301]<=26'd23456209;
ROM1[5302]<=26'd1976022; ROM2[5302]<=26'd11175952; ROM3[5302]<=26'd9745473; ROM4[5302]<=26'd23458160;
ROM1[5303]<=26'd1974188; ROM2[5303]<=26'd11178155; ROM3[5303]<=26'd9751379; ROM4[5303]<=26'd23461557;
ROM1[5304]<=26'd1972126; ROM2[5304]<=26'd11181229; ROM3[5304]<=26'd9754432; ROM4[5304]<=26'd23465379;
ROM1[5305]<=26'd1974030; ROM2[5305]<=26'd11181847; ROM3[5305]<=26'd9754032; ROM4[5305]<=26'd23465202;
ROM1[5306]<=26'd1977758; ROM2[5306]<=26'd11178842; ROM3[5306]<=26'd9746997; ROM4[5306]<=26'd23461206;
ROM1[5307]<=26'd1986565; ROM2[5307]<=26'd11177150; ROM3[5307]<=26'd9740033; ROM4[5307]<=26'd23458139;
ROM1[5308]<=26'd1987611; ROM2[5308]<=26'd11175140; ROM3[5308]<=26'd9736466; ROM4[5308]<=26'd23455768;
ROM1[5309]<=26'd1982794; ROM2[5309]<=26'd11174366; ROM3[5309]<=26'd9738909; ROM4[5309]<=26'd23456589;
ROM1[5310]<=26'd1978154; ROM2[5310]<=26'd11174734; ROM3[5310]<=26'd9745080; ROM4[5310]<=26'd23458601;
ROM1[5311]<=26'd1974574; ROM2[5311]<=26'd11173686; ROM3[5311]<=26'd9747806; ROM4[5311]<=26'd23458700;
ROM1[5312]<=26'd1969597; ROM2[5312]<=26'd11177038; ROM3[5312]<=26'd9753220; ROM4[5312]<=26'd23461314;
ROM1[5313]<=26'd1967299; ROM2[5313]<=26'd11177819; ROM3[5313]<=26'd9752556; ROM4[5313]<=26'd23460160;
ROM1[5314]<=26'd1975879; ROM2[5314]<=26'd11177659; ROM3[5314]<=26'd9748462; ROM4[5314]<=26'd23459424;
ROM1[5315]<=26'd1984169; ROM2[5315]<=26'd11177571; ROM3[5315]<=26'd9740698; ROM4[5315]<=26'd23456477;
ROM1[5316]<=26'd1986550; ROM2[5316]<=26'd11173424; ROM3[5316]<=26'd9735220; ROM4[5316]<=26'd23453046;
ROM1[5317]<=26'd1985454; ROM2[5317]<=26'd11173827; ROM3[5317]<=26'd9739905; ROM4[5317]<=26'd23454821;
ROM1[5318]<=26'd1979635; ROM2[5318]<=26'd11175639; ROM3[5318]<=26'd9744633; ROM4[5318]<=26'd23456068;
ROM1[5319]<=26'd1978024; ROM2[5319]<=26'd11177782; ROM3[5319]<=26'd9751441; ROM4[5319]<=26'd23460389;
ROM1[5320]<=26'd1973342; ROM2[5320]<=26'd11175502; ROM3[5320]<=26'd9754033; ROM4[5320]<=26'd23461048;
ROM1[5321]<=26'd1967327; ROM2[5321]<=26'd11170624; ROM3[5321]<=26'd9751482; ROM4[5321]<=26'd23457104;
ROM1[5322]<=26'd1975333; ROM2[5322]<=26'd11176903; ROM3[5322]<=26'd9754980; ROM4[5322]<=26'd23462064;
ROM1[5323]<=26'd1987331; ROM2[5323]<=26'd11179278; ROM3[5323]<=26'd9750036; ROM4[5323]<=26'd23460686;
ROM1[5324]<=26'd1991221; ROM2[5324]<=26'd11175949; ROM3[5324]<=26'd9738344; ROM4[5324]<=26'd23452615;
ROM1[5325]<=26'd1991293; ROM2[5325]<=26'd11180288; ROM3[5325]<=26'd9738053; ROM4[5325]<=26'd23453240;
ROM1[5326]<=26'd1976404; ROM2[5326]<=26'd11171049; ROM3[5326]<=26'd9731666; ROM4[5326]<=26'd23444926;
ROM1[5327]<=26'd1965502; ROM2[5327]<=26'd11164771; ROM3[5327]<=26'd9731316; ROM4[5327]<=26'd23440913;
ROM1[5328]<=26'd1965612; ROM2[5328]<=26'd11170084; ROM3[5328]<=26'd9739218; ROM4[5328]<=26'd23447992;
ROM1[5329]<=26'd1962165; ROM2[5329]<=26'd11171186; ROM3[5329]<=26'd9740061; ROM4[5329]<=26'd23448274;
ROM1[5330]<=26'd1967850; ROM2[5330]<=26'd11176083; ROM3[5330]<=26'd9740369; ROM4[5330]<=26'd23449262;
ROM1[5331]<=26'd1980087; ROM2[5331]<=26'd11181652; ROM3[5331]<=26'd9738489; ROM4[5331]<=26'd23453469;
ROM1[5332]<=26'd1988364; ROM2[5332]<=26'd11177962; ROM3[5332]<=26'd9731079; ROM4[5332]<=26'd23450134;
ROM1[5333]<=26'd1990153; ROM2[5333]<=26'd11177320; ROM3[5333]<=26'd9731398; ROM4[5333]<=26'd23450989;
ROM1[5334]<=26'd1984787; ROM2[5334]<=26'd11177064; ROM3[5334]<=26'd9734527; ROM4[5334]<=26'd23451487;
ROM1[5335]<=26'd1977966; ROM2[5335]<=26'd11173905; ROM3[5335]<=26'd9736423; ROM4[5335]<=26'd23450218;
ROM1[5336]<=26'd1977537; ROM2[5336]<=26'd11178462; ROM3[5336]<=26'd9743586; ROM4[5336]<=26'd23454700;
ROM1[5337]<=26'd1971984; ROM2[5337]<=26'd11177604; ROM3[5337]<=26'd9746829; ROM4[5337]<=26'd23455789;
ROM1[5338]<=26'd1970955; ROM2[5338]<=26'd11176699; ROM3[5338]<=26'd9746599; ROM4[5338]<=26'd23457400;
ROM1[5339]<=26'd1981395; ROM2[5339]<=26'd11179470; ROM3[5339]<=26'd9746771; ROM4[5339]<=26'd23459103;
ROM1[5340]<=26'd1992793; ROM2[5340]<=26'd11177474; ROM3[5340]<=26'd9741040; ROM4[5340]<=26'd23456496;
ROM1[5341]<=26'd1998557; ROM2[5341]<=26'd11177997; ROM3[5341]<=26'd9740028; ROM4[5341]<=26'd23458846;
ROM1[5342]<=26'd1994246; ROM2[5342]<=26'd11177031; ROM3[5342]<=26'd9742361; ROM4[5342]<=26'd23460760;
ROM1[5343]<=26'd1983583; ROM2[5343]<=26'd11172770; ROM3[5343]<=26'd9743191; ROM4[5343]<=26'd23458176;
ROM1[5344]<=26'd1979953; ROM2[5344]<=26'd11173569; ROM3[5344]<=26'd9748125; ROM4[5344]<=26'd23460056;
ROM1[5345]<=26'd1975026; ROM2[5345]<=26'd11173378; ROM3[5345]<=26'd9751129; ROM4[5345]<=26'd23459491;
ROM1[5346]<=26'd1971720; ROM2[5346]<=26'd11172509; ROM3[5346]<=26'd9750837; ROM4[5346]<=26'd23458270;
ROM1[5347]<=26'd1977349; ROM2[5347]<=26'd11175485; ROM3[5347]<=26'd9748608; ROM4[5347]<=26'd23459494;
ROM1[5348]<=26'd1991636; ROM2[5348]<=26'd11177488; ROM3[5348]<=26'd9745347; ROM4[5348]<=26'd23461179;
ROM1[5349]<=26'd2001762; ROM2[5349]<=26'd11177667; ROM3[5349]<=26'd9743675; ROM4[5349]<=26'd23463365;
ROM1[5350]<=26'd1999259; ROM2[5350]<=26'd11177121; ROM3[5350]<=26'd9746126; ROM4[5350]<=26'd23463018;
ROM1[5351]<=26'd1991656; ROM2[5351]<=26'd11175154; ROM3[5351]<=26'd9747639; ROM4[5351]<=26'd23462759;
ROM1[5352]<=26'd1981764; ROM2[5352]<=26'd11172656; ROM3[5352]<=26'd9749259; ROM4[5352]<=26'd23461797;
ROM1[5353]<=26'd1978578; ROM2[5353]<=26'd11175319; ROM3[5353]<=26'd9753725; ROM4[5353]<=26'd23464915;
ROM1[5354]<=26'd1979097; ROM2[5354]<=26'd11180723; ROM3[5354]<=26'd9756359; ROM4[5354]<=26'd23468253;
ROM1[5355]<=26'd1981629; ROM2[5355]<=26'd11181535; ROM3[5355]<=26'd9756284; ROM4[5355]<=26'd23468013;
ROM1[5356]<=26'd1987725; ROM2[5356]<=26'd11180131; ROM3[5356]<=26'd9750396; ROM4[5356]<=26'd23465397;
ROM1[5357]<=26'd1998457; ROM2[5357]<=26'd11179907; ROM3[5357]<=26'd9742693; ROM4[5357]<=26'd23464405;
ROM1[5358]<=26'd1999083; ROM2[5358]<=26'd11177584; ROM3[5358]<=26'd9741286; ROM4[5358]<=26'd23463389;
ROM1[5359]<=26'd1988192; ROM2[5359]<=26'd11173527; ROM3[5359]<=26'd9741141; ROM4[5359]<=26'd23461365;
ROM1[5360]<=26'd1979599; ROM2[5360]<=26'd11171040; ROM3[5360]<=26'd9741907; ROM4[5360]<=26'd23460608;
ROM1[5361]<=26'd1973965; ROM2[5361]<=26'd11168821; ROM3[5361]<=26'd9742582; ROM4[5361]<=26'd23458920;
ROM1[5362]<=26'd1965799; ROM2[5362]<=26'd11165186; ROM3[5362]<=26'd9742587; ROM4[5362]<=26'd23456001;
ROM1[5363]<=26'd1966298; ROM2[5363]<=26'd11165095; ROM3[5363]<=26'd9743118; ROM4[5363]<=26'd23454826;
ROM1[5364]<=26'd1976737; ROM2[5364]<=26'd11171725; ROM3[5364]<=26'd9745168; ROM4[5364]<=26'd23458725;
ROM1[5365]<=26'd1993033; ROM2[5365]<=26'd11179963; ROM3[5365]<=26'd9747106; ROM4[5365]<=26'd23465519;
ROM1[5366]<=26'd1993447; ROM2[5366]<=26'd11172631; ROM3[5366]<=26'd9737644; ROM4[5366]<=26'd23459207;
ROM1[5367]<=26'd1983162; ROM2[5367]<=26'd11164495; ROM3[5367]<=26'd9733578; ROM4[5367]<=26'd23452616;
ROM1[5368]<=26'd1980428; ROM2[5368]<=26'd11167065; ROM3[5368]<=26'd9740499; ROM4[5368]<=26'd23456807;
ROM1[5369]<=26'd1972714; ROM2[5369]<=26'd11164557; ROM3[5369]<=26'd9741396; ROM4[5369]<=26'd23454917;
ROM1[5370]<=26'd1967638; ROM2[5370]<=26'd11166352; ROM3[5370]<=26'd9747018; ROM4[5370]<=26'd23458098;
ROM1[5371]<=26'd1969263; ROM2[5371]<=26'd11171706; ROM3[5371]<=26'd9752949; ROM4[5371]<=26'd23462835;
ROM1[5372]<=26'd1975967; ROM2[5372]<=26'd11173161; ROM3[5372]<=26'd9752161; ROM4[5372]<=26'd23464315;
ROM1[5373]<=26'd1987106; ROM2[5373]<=26'd11172214; ROM3[5373]<=26'd9744793; ROM4[5373]<=26'd23461430;
ROM1[5374]<=26'd1990542; ROM2[5374]<=26'd11168187; ROM3[5374]<=26'd9734878; ROM4[5374]<=26'd23454824;
ROM1[5375]<=26'd1990706; ROM2[5375]<=26'd11171098; ROM3[5375]<=26'd9736134; ROM4[5375]<=26'd23455759;
ROM1[5376]<=26'd1983966; ROM2[5376]<=26'd11170354; ROM3[5376]<=26'd9740102; ROM4[5376]<=26'd23455722;
ROM1[5377]<=26'd1976713; ROM2[5377]<=26'd11168683; ROM3[5377]<=26'd9742778; ROM4[5377]<=26'd23456538;
ROM1[5378]<=26'd1974646; ROM2[5378]<=26'd11172082; ROM3[5378]<=26'd9747607; ROM4[5378]<=26'd23459666;
ROM1[5379]<=26'd1966529; ROM2[5379]<=26'd11168426; ROM3[5379]<=26'd9746040; ROM4[5379]<=26'd23456347;
ROM1[5380]<=26'd1964825; ROM2[5380]<=26'd11165400; ROM3[5380]<=26'd9741148; ROM4[5380]<=26'd23451379;
ROM1[5381]<=26'd1974611; ROM2[5381]<=26'd11166576; ROM3[5381]<=26'd9736954; ROM4[5381]<=26'd23448285;
ROM1[5382]<=26'd1990607; ROM2[5382]<=26'd11170853; ROM3[5382]<=26'd9735583; ROM4[5382]<=26'd23452355;
ROM1[5383]<=26'd1992583; ROM2[5383]<=26'd11171390; ROM3[5383]<=26'd9736526; ROM4[5383]<=26'd23455053;
ROM1[5384]<=26'd1988043; ROM2[5384]<=26'd11172893; ROM3[5384]<=26'd9741337; ROM4[5384]<=26'd23456753;
ROM1[5385]<=26'd1979566; ROM2[5385]<=26'd11171147; ROM3[5385]<=26'd9744122; ROM4[5385]<=26'd23455678;
ROM1[5386]<=26'd1973277; ROM2[5386]<=26'd11169146; ROM3[5386]<=26'd9745328; ROM4[5386]<=26'd23454000;
ROM1[5387]<=26'd1970724; ROM2[5387]<=26'd11168724; ROM3[5387]<=26'd9748161; ROM4[5387]<=26'd23453716;
ROM1[5388]<=26'd1968708; ROM2[5388]<=26'd11167570; ROM3[5388]<=26'd9746218; ROM4[5388]<=26'd23451086;
ROM1[5389]<=26'd1973903; ROM2[5389]<=26'd11167184; ROM3[5389]<=26'd9743123; ROM4[5389]<=26'd23450469;
ROM1[5390]<=26'd1988321; ROM2[5390]<=26'd11169287; ROM3[5390]<=26'd9741165; ROM4[5390]<=26'd23452355;
ROM1[5391]<=26'd1997688; ROM2[5391]<=26'd11171879; ROM3[5391]<=26'd9739567; ROM4[5391]<=26'd23454089;
ROM1[5392]<=26'd1988648; ROM2[5392]<=26'd11165029; ROM3[5392]<=26'd9735228; ROM4[5392]<=26'd23449330;
ROM1[5393]<=26'd1982788; ROM2[5393]<=26'd11165556; ROM3[5393]<=26'd9740657; ROM4[5393]<=26'd23451066;
ROM1[5394]<=26'd1978959; ROM2[5394]<=26'd11168060; ROM3[5394]<=26'd9744650; ROM4[5394]<=26'd23453512;
ROM1[5395]<=26'd1971889; ROM2[5395]<=26'd11169065; ROM3[5395]<=26'd9748688; ROM4[5395]<=26'd23455485;
ROM1[5396]<=26'd1974189; ROM2[5396]<=26'd11174014; ROM3[5396]<=26'd9753585; ROM4[5396]<=26'd23458942;
ROM1[5397]<=26'd1979809; ROM2[5397]<=26'd11174160; ROM3[5397]<=26'd9751457; ROM4[5397]<=26'd23457560;
ROM1[5398]<=26'd1988864; ROM2[5398]<=26'd11171515; ROM3[5398]<=26'd9744068; ROM4[5398]<=26'd23453812;
ROM1[5399]<=26'd1995354; ROM2[5399]<=26'd11169151; ROM3[5399]<=26'd9736424; ROM4[5399]<=26'd23450708;
ROM1[5400]<=26'd1992058; ROM2[5400]<=26'd11167047; ROM3[5400]<=26'd9737336; ROM4[5400]<=26'd23451347;
ROM1[5401]<=26'd1988346; ROM2[5401]<=26'd11168861; ROM3[5401]<=26'd9743030; ROM4[5401]<=26'd23453825;
ROM1[5402]<=26'd1984399; ROM2[5402]<=26'd11172452; ROM3[5402]<=26'd9750598; ROM4[5402]<=26'd23457179;
ROM1[5403]<=26'd1979682; ROM2[5403]<=26'd11172567; ROM3[5403]<=26'd9755412; ROM4[5403]<=26'd23459803;
ROM1[5404]<=26'd1975324; ROM2[5404]<=26'd11170994; ROM3[5404]<=26'd9756346; ROM4[5404]<=26'd23461038;
ROM1[5405]<=26'd1976258; ROM2[5405]<=26'd11168579; ROM3[5405]<=26'd9754549; ROM4[5405]<=26'd23459707;
ROM1[5406]<=26'd1987370; ROM2[5406]<=26'd11169753; ROM3[5406]<=26'd9748525; ROM4[5406]<=26'd23458981;
ROM1[5407]<=26'd1996489; ROM2[5407]<=26'd11170071; ROM3[5407]<=26'd9738838; ROM4[5407]<=26'd23455846;
ROM1[5408]<=26'd1999227; ROM2[5408]<=26'd11171401; ROM3[5408]<=26'd9739439; ROM4[5408]<=26'd23456139;
ROM1[5409]<=26'd1998929; ROM2[5409]<=26'd11176970; ROM3[5409]<=26'd9747061; ROM4[5409]<=26'd23462447;
ROM1[5410]<=26'd1996018; ROM2[5410]<=26'd11180975; ROM3[5410]<=26'd9756760; ROM4[5410]<=26'd23467742;
ROM1[5411]<=26'd1985755; ROM2[5411]<=26'd11172787; ROM3[5411]<=26'd9754650; ROM4[5411]<=26'd23462683;
ROM1[5412]<=26'd1972383; ROM2[5412]<=26'd11165031; ROM3[5412]<=26'd9749467; ROM4[5412]<=26'd23455378;
ROM1[5413]<=26'd1970219; ROM2[5413]<=26'd11161782; ROM3[5413]<=26'd9745996; ROM4[5413]<=26'd23452224;
ROM1[5414]<=26'd1976334; ROM2[5414]<=26'd11159761; ROM3[5414]<=26'd9739312; ROM4[5414]<=26'd23449845;
ROM1[5415]<=26'd1992635; ROM2[5415]<=26'd11164734; ROM3[5415]<=26'd9738632; ROM4[5415]<=26'd23452121;
ROM1[5416]<=26'd1999405; ROM2[5416]<=26'd11168514; ROM3[5416]<=26'd9738093; ROM4[5416]<=26'd23454189;
ROM1[5417]<=26'd1998630; ROM2[5417]<=26'd11173353; ROM3[5417]<=26'd9743028; ROM4[5417]<=26'd23459437;
ROM1[5418]<=26'd1983968; ROM2[5418]<=26'd11163944; ROM3[5418]<=26'd9739402; ROM4[5418]<=26'd23452113;
ROM1[5419]<=26'd1971870; ROM2[5419]<=26'd11157532; ROM3[5419]<=26'd9735694; ROM4[5419]<=26'd23445768;
ROM1[5420]<=26'd1969796; ROM2[5420]<=26'd11161506; ROM3[5420]<=26'd9740155; ROM4[5420]<=26'd23450283;
ROM1[5421]<=26'd1963531; ROM2[5421]<=26'd11157379; ROM3[5421]<=26'd9736727; ROM4[5421]<=26'd23446682;
ROM1[5422]<=26'd1967625; ROM2[5422]<=26'd11157111; ROM3[5422]<=26'd9733234; ROM4[5422]<=26'd23445248;
ROM1[5423]<=26'd1988576; ROM2[5423]<=26'd11167346; ROM3[5423]<=26'd9734527; ROM4[5423]<=26'd23453374;
ROM1[5424]<=26'd2004990; ROM2[5424]<=26'd11172422; ROM3[5424]<=26'd9736751; ROM4[5424]<=26'd23458541;
ROM1[5425]<=26'd2005762; ROM2[5425]<=26'd11173836; ROM3[5425]<=26'd9740406; ROM4[5425]<=26'd23461866;
ROM1[5426]<=26'd2003603; ROM2[5426]<=26'd11181515; ROM3[5426]<=26'd9749394; ROM4[5426]<=26'd23469219;
ROM1[5427]<=26'd1995251; ROM2[5427]<=26'd11181312; ROM3[5427]<=26'd9755119; ROM4[5427]<=26'd23469607;
ROM1[5428]<=26'd1987725; ROM2[5428]<=26'd11178564; ROM3[5428]<=26'd9755809; ROM4[5428]<=26'd23467701;
ROM1[5429]<=26'd1983942; ROM2[5429]<=26'd11178014; ROM3[5429]<=26'd9756910; ROM4[5429]<=26'd23467698;
ROM1[5430]<=26'd1978165; ROM2[5430]<=26'd11169728; ROM3[5430]<=26'd9749378; ROM4[5430]<=26'd23459133;
ROM1[5431]<=26'd1990096; ROM2[5431]<=26'd11169155; ROM3[5431]<=26'd9743539; ROM4[5431]<=26'd23458433;
ROM1[5432]<=26'd2005393; ROM2[5432]<=26'd11172431; ROM3[5432]<=26'd9740785; ROM4[5432]<=26'd23460422;
ROM1[5433]<=26'd2003571; ROM2[5433]<=26'd11170805; ROM3[5433]<=26'd9738620; ROM4[5433]<=26'd23457560;
ROM1[5434]<=26'd1999570; ROM2[5434]<=26'd11171499; ROM3[5434]<=26'd9744299; ROM4[5434]<=26'd23461279;
ROM1[5435]<=26'd1989296; ROM2[5435]<=26'd11169959; ROM3[5435]<=26'd9746220; ROM4[5435]<=26'd23460216;
ROM1[5436]<=26'd1980875; ROM2[5436]<=26'd11167538; ROM3[5436]<=26'd9745101; ROM4[5436]<=26'd23458123;
ROM1[5437]<=26'd1972664; ROM2[5437]<=26'd11163579; ROM3[5437]<=26'd9743371; ROM4[5437]<=26'd23453248;
ROM1[5438]<=26'd1975847; ROM2[5438]<=26'd11166083; ROM3[5438]<=26'd9742615; ROM4[5438]<=26'd23452328;
ROM1[5439]<=26'd1986320; ROM2[5439]<=26'd11167927; ROM3[5439]<=26'd9742093; ROM4[5439]<=26'd23453187;
ROM1[5440]<=26'd1997194; ROM2[5440]<=26'd11168945; ROM3[5440]<=26'd9737907; ROM4[5440]<=26'd23452707;
ROM1[5441]<=26'd2004580; ROM2[5441]<=26'd11173075; ROM3[5441]<=26'd9735789; ROM4[5441]<=26'd23454994;
ROM1[5442]<=26'd2003190; ROM2[5442]<=26'd11175749; ROM3[5442]<=26'd9737553; ROM4[5442]<=26'd23457139;
ROM1[5443]<=26'd1993402; ROM2[5443]<=26'd11172597; ROM3[5443]<=26'd9738407; ROM4[5443]<=26'd23455781;
ROM1[5444]<=26'd1986078; ROM2[5444]<=26'd11169554; ROM3[5444]<=26'd9739763; ROM4[5444]<=26'd23452806;
ROM1[5445]<=26'd1983299; ROM2[5445]<=26'd11170693; ROM3[5445]<=26'd9744694; ROM4[5445]<=26'd23455085;
ROM1[5446]<=26'd1984464; ROM2[5446]<=26'd11174792; ROM3[5446]<=26'd9749724; ROM4[5446]<=26'd23459912;
ROM1[5447]<=26'd1991000; ROM2[5447]<=26'd11176798; ROM3[5447]<=26'd9749768; ROM4[5447]<=26'd23460656;
ROM1[5448]<=26'd2002925; ROM2[5448]<=26'd11174902; ROM3[5448]<=26'd9744592; ROM4[5448]<=26'd23460300;
ROM1[5449]<=26'd2010184; ROM2[5449]<=26'd11172914; ROM3[5449]<=26'd9739798; ROM4[5449]<=26'd23458850;
ROM1[5450]<=26'd2003591; ROM2[5450]<=26'd11168393; ROM3[5450]<=26'd9737426; ROM4[5450]<=26'd23454787;
ROM1[5451]<=26'd1997899; ROM2[5451]<=26'd11167538; ROM3[5451]<=26'd9739509; ROM4[5451]<=26'd23455733;
ROM1[5452]<=26'd1991813; ROM2[5452]<=26'd11167624; ROM3[5452]<=26'd9741048; ROM4[5452]<=26'd23455077;
ROM1[5453]<=26'd1982296; ROM2[5453]<=26'd11163429; ROM3[5453]<=26'd9740991; ROM4[5453]<=26'd23452088;
ROM1[5454]<=26'd1976949; ROM2[5454]<=26'd11160933; ROM3[5454]<=26'd9742615; ROM4[5454]<=26'd23453058;
ROM1[5455]<=26'd1980964; ROM2[5455]<=26'd11162232; ROM3[5455]<=26'd9744133; ROM4[5455]<=26'd23453958;
ROM1[5456]<=26'd1989837; ROM2[5456]<=26'd11162748; ROM3[5456]<=26'd9739896; ROM4[5456]<=26'd23450010;
ROM1[5457]<=26'd2000329; ROM2[5457]<=26'd11162576; ROM3[5457]<=26'd9732725; ROM4[5457]<=26'd23448242;
ROM1[5458]<=26'd2010042; ROM2[5458]<=26'd11171070; ROM3[5458]<=26'd9739355; ROM4[5458]<=26'd23456558;
ROM1[5459]<=26'd2004211; ROM2[5459]<=26'd11171190; ROM3[5459]<=26'd9742619; ROM4[5459]<=26'd23457120;
ROM1[5460]<=26'd1992519; ROM2[5460]<=26'd11165687; ROM3[5460]<=26'd9741688; ROM4[5460]<=26'd23453917;
ROM1[5461]<=26'd1994224; ROM2[5461]<=26'd11170651; ROM3[5461]<=26'd9749573; ROM4[5461]<=26'd23459922;
ROM1[5462]<=26'd1989225; ROM2[5462]<=26'd11170146; ROM3[5462]<=26'd9751206; ROM4[5462]<=26'd23459209;
ROM1[5463]<=26'd1988416; ROM2[5463]<=26'd11170170; ROM3[5463]<=26'd9749082; ROM4[5463]<=26'd23458107;
ROM1[5464]<=26'd1997882; ROM2[5464]<=26'd11172851; ROM3[5464]<=26'd9747672; ROM4[5464]<=26'd23458515;
ROM1[5465]<=26'd2005936; ROM2[5465]<=26'd11171438; ROM3[5465]<=26'd9738251; ROM4[5465]<=26'd23454472;
ROM1[5466]<=26'd2005000; ROM2[5466]<=26'd11165087; ROM3[5466]<=26'd9730288; ROM4[5466]<=26'd23448220;
ROM1[5467]<=26'd1999047; ROM2[5467]<=26'd11163448; ROM3[5467]<=26'd9732514; ROM4[5467]<=26'd23448875;
ROM1[5468]<=26'd1995907; ROM2[5468]<=26'd11165487; ROM3[5468]<=26'd9739382; ROM4[5468]<=26'd23455000;
ROM1[5469]<=26'd1997924; ROM2[5469]<=26'd11169406; ROM3[5469]<=26'd9748115; ROM4[5469]<=26'd23459691;
ROM1[5470]<=26'd2002297; ROM2[5470]<=26'd11176498; ROM3[5470]<=26'd9758826; ROM4[5470]<=26'd23466923;
ROM1[5471]<=26'd1994268; ROM2[5471]<=26'd11169086; ROM3[5471]<=26'd9752255; ROM4[5471]<=26'd23458942;
ROM1[5472]<=26'd1990307; ROM2[5472]<=26'd11161167; ROM3[5472]<=26'd9744146; ROM4[5472]<=26'd23451829;
ROM1[5473]<=26'd2002666; ROM2[5473]<=26'd11162816; ROM3[5473]<=26'd9741144; ROM4[5473]<=26'd23453333;
ROM1[5474]<=26'd2006265; ROM2[5474]<=26'd11158972; ROM3[5474]<=26'd9732787; ROM4[5474]<=26'd23447923;
ROM1[5475]<=26'd2006857; ROM2[5475]<=26'd11162123; ROM3[5475]<=26'd9737996; ROM4[5475]<=26'd23451774;
ROM1[5476]<=26'd2003219; ROM2[5476]<=26'd11163116; ROM3[5476]<=26'd9740210; ROM4[5476]<=26'd23452176;
ROM1[5477]<=26'd1991965; ROM2[5477]<=26'd11156616; ROM3[5477]<=26'd9737418; ROM4[5477]<=26'd23446199;
ROM1[5478]<=26'd1982422; ROM2[5478]<=26'd11152299; ROM3[5478]<=26'd9737127; ROM4[5478]<=26'd23443902;
ROM1[5479]<=26'd1978074; ROM2[5479]<=26'd11151496; ROM3[5479]<=26'd9739212; ROM4[5479]<=26'd23443984;
ROM1[5480]<=26'd1984121; ROM2[5480]<=26'd11155958; ROM3[5480]<=26'd9742878; ROM4[5480]<=26'd23447168;
ROM1[5481]<=26'd1996841; ROM2[5481]<=26'd11159641; ROM3[5481]<=26'd9741112; ROM4[5481]<=26'd23449262;
ROM1[5482]<=26'd2010709; ROM2[5482]<=26'd11163057; ROM3[5482]<=26'd9736959; ROM4[5482]<=26'd23451056;
ROM1[5483]<=26'd2008210; ROM2[5483]<=26'd11162753; ROM3[5483]<=26'd9733391; ROM4[5483]<=26'd23449832;
ROM1[5484]<=26'd1999972; ROM2[5484]<=26'd11162096; ROM3[5484]<=26'd9735197; ROM4[5484]<=26'd23449758;
ROM1[5485]<=26'd1992428; ROM2[5485]<=26'd11161711; ROM3[5485]<=26'd9737912; ROM4[5485]<=26'd23449464;
ROM1[5486]<=26'd1985177; ROM2[5486]<=26'd11158988; ROM3[5486]<=26'd9737404; ROM4[5486]<=26'd23447107;
ROM1[5487]<=26'd1985872; ROM2[5487]<=26'd11162495; ROM3[5487]<=26'd9743018; ROM4[5487]<=26'd23451415;
ROM1[5488]<=26'd1991486; ROM2[5488]<=26'd11169099; ROM3[5488]<=26'd9748162; ROM4[5488]<=26'd23457688;
ROM1[5489]<=26'd1995989; ROM2[5489]<=26'd11166482; ROM3[5489]<=26'd9743130; ROM4[5489]<=26'd23455440;
ROM1[5490]<=26'd2005889; ROM2[5490]<=26'd11164171; ROM3[5490]<=26'd9735320; ROM4[5490]<=26'd23451032;
ROM1[5491]<=26'd2010377; ROM2[5491]<=26'd11163731; ROM3[5491]<=26'd9732957; ROM4[5491]<=26'd23451288;
ROM1[5492]<=26'd2003733; ROM2[5492]<=26'd11160515; ROM3[5492]<=26'd9732659; ROM4[5492]<=26'd23449408;
ROM1[5493]<=26'd1993779; ROM2[5493]<=26'd11157967; ROM3[5493]<=26'd9733344; ROM4[5493]<=26'd23446896;
ROM1[5494]<=26'd1990564; ROM2[5494]<=26'd11158390; ROM3[5494]<=26'd9737676; ROM4[5494]<=26'd23449168;
ROM1[5495]<=26'd1987642; ROM2[5495]<=26'd11160827; ROM3[5495]<=26'd9743576; ROM4[5495]<=26'd23452566;
ROM1[5496]<=26'd1985201; ROM2[5496]<=26'd11160139; ROM3[5496]<=26'd9742914; ROM4[5496]<=26'd23451762;
ROM1[5497]<=26'd1990061; ROM2[5497]<=26'd11158669; ROM3[5497]<=26'd9740461; ROM4[5497]<=26'd23450681;
ROM1[5498]<=26'd2001591; ROM2[5498]<=26'd11159894; ROM3[5498]<=26'd9737705; ROM4[5498]<=26'd23451795;
ROM1[5499]<=26'd2013546; ROM2[5499]<=26'd11163576; ROM3[5499]<=26'd9735598; ROM4[5499]<=26'd23453549;
ROM1[5500]<=26'd2011756; ROM2[5500]<=26'd11162898; ROM3[5500]<=26'd9736280; ROM4[5500]<=26'd23452615;
ROM1[5501]<=26'd2011572; ROM2[5501]<=26'd11167738; ROM3[5501]<=26'd9742930; ROM4[5501]<=26'd23457235;
ROM1[5502]<=26'd2015883; ROM2[5502]<=26'd11176601; ROM3[5502]<=26'd9755285; ROM4[5502]<=26'd23466776;
ROM1[5503]<=26'd2005323; ROM2[5503]<=26'd11169951; ROM3[5503]<=26'd9751785; ROM4[5503]<=26'd23459536;
ROM1[5504]<=26'd1999422; ROM2[5504]<=26'd11167917; ROM3[5504]<=26'd9749527; ROM4[5504]<=26'd23456589;
ROM1[5505]<=26'd1999690; ROM2[5505]<=26'd11166086; ROM3[5505]<=26'd9746372; ROM4[5505]<=26'd23453662;
ROM1[5506]<=26'd2001012; ROM2[5506]<=26'd11157678; ROM3[5506]<=26'd9732722; ROM4[5506]<=26'd23441928;
ROM1[5507]<=26'd2015348; ROM2[5507]<=26'd11160431; ROM3[5507]<=26'd9729901; ROM4[5507]<=26'd23444287;
ROM1[5508]<=26'd2017661; ROM2[5508]<=26'd11163220; ROM3[5508]<=26'd9733620; ROM4[5508]<=26'd23446560;
ROM1[5509]<=26'd2009224; ROM2[5509]<=26'd11162265; ROM3[5509]<=26'd9735112; ROM4[5509]<=26'd23444047;
ROM1[5510]<=26'd1998235; ROM2[5510]<=26'd11158402; ROM3[5510]<=26'd9735897; ROM4[5510]<=26'd23441645;
ROM1[5511]<=26'd1988513; ROM2[5511]<=26'd11154904; ROM3[5511]<=26'd9735477; ROM4[5511]<=26'd23439464;
ROM1[5512]<=26'd1982119; ROM2[5512]<=26'd11153025; ROM3[5512]<=26'd9733667; ROM4[5512]<=26'd23437754;
ROM1[5513]<=26'd1980996; ROM2[5513]<=26'd11150255; ROM3[5513]<=26'd9731618; ROM4[5513]<=26'd23436003;
ROM1[5514]<=26'd1992885; ROM2[5514]<=26'd11158685; ROM3[5514]<=26'd9732963; ROM4[5514]<=26'd23441381;
ROM1[5515]<=26'd2020212; ROM2[5515]<=26'd11174064; ROM3[5515]<=26'd9739220; ROM4[5515]<=26'd23452936;
ROM1[5516]<=26'd2019429; ROM2[5516]<=26'd11166740; ROM3[5516]<=26'd9731843; ROM4[5516]<=26'd23448286;
ROM1[5517]<=26'd2003302; ROM2[5517]<=26'd11156386; ROM3[5517]<=26'd9725126; ROM4[5517]<=26'd23441614;
ROM1[5518]<=26'd2000721; ROM2[5518]<=26'd11159939; ROM3[5518]<=26'd9731693; ROM4[5518]<=26'd23446675;
ROM1[5519]<=26'd1993523; ROM2[5519]<=26'd11157948; ROM3[5519]<=26'd9732897; ROM4[5519]<=26'd23445392;
ROM1[5520]<=26'd1987828; ROM2[5520]<=26'd11157020; ROM3[5520]<=26'd9733498; ROM4[5520]<=26'd23444977;
ROM1[5521]<=26'd1985415; ROM2[5521]<=26'd11157920; ROM3[5521]<=26'd9734406; ROM4[5521]<=26'd23445328;
ROM1[5522]<=26'd1987232; ROM2[5522]<=26'd11153995; ROM3[5522]<=26'd9729393; ROM4[5522]<=26'd23441519;
ROM1[5523]<=26'd1996420; ROM2[5523]<=26'd11151684; ROM3[5523]<=26'd9721330; ROM4[5523]<=26'd23438864;
ROM1[5524]<=26'd2012784; ROM2[5524]<=26'd11158539; ROM3[5524]<=26'd9725311; ROM4[5524]<=26'd23445633;
ROM1[5525]<=26'd2018349; ROM2[5525]<=26'd11166104; ROM3[5525]<=26'd9732886; ROM4[5525]<=26'd23452113;
ROM1[5526]<=26'd2006779; ROM2[5526]<=26'd11162164; ROM3[5526]<=26'd9732926; ROM4[5526]<=26'd23448143;
ROM1[5527]<=26'd1998083; ROM2[5527]<=26'd11157239; ROM3[5527]<=26'd9733896; ROM4[5527]<=26'd23445360;
ROM1[5528]<=26'd1994453; ROM2[5528]<=26'd11159331; ROM3[5528]<=26'd9738958; ROM4[5528]<=26'd23448858;
ROM1[5529]<=26'd1991640; ROM2[5529]<=26'd11160965; ROM3[5529]<=26'd9745407; ROM4[5529]<=26'd23452587;
ROM1[5530]<=26'd1998193; ROM2[5530]<=26'd11164131; ROM3[5530]<=26'd9749982; ROM4[5530]<=26'd23457482;
ROM1[5531]<=26'd2011036; ROM2[5531]<=26'd11166849; ROM3[5531]<=26'd9749008; ROM4[5531]<=26'd23459320;
ROM1[5532]<=26'd2022946; ROM2[5532]<=26'd11166743; ROM3[5532]<=26'd9745011; ROM4[5532]<=26'd23457653;
ROM1[5533]<=26'd2026193; ROM2[5533]<=26'd11167558; ROM3[5533]<=26'd9747498; ROM4[5533]<=26'd23459738;
ROM1[5534]<=26'd2017597; ROM2[5534]<=26'd11163788; ROM3[5534]<=26'd9746557; ROM4[5534]<=26'd23455783;
ROM1[5535]<=26'd2013709; ROM2[5535]<=26'd11166852; ROM3[5535]<=26'd9751044; ROM4[5535]<=26'd23457839;
ROM1[5536]<=26'd2014054; ROM2[5536]<=26'd11173951; ROM3[5536]<=26'd9759034; ROM4[5536]<=26'd23463367;
ROM1[5537]<=26'd2001585; ROM2[5537]<=26'd11167360; ROM3[5537]<=26'd9754593; ROM4[5537]<=26'd23455846;
ROM1[5538]<=26'd1992750; ROM2[5538]<=26'd11158417; ROM3[5538]<=26'd9744910; ROM4[5538]<=26'd23447656;
ROM1[5539]<=26'd1996895; ROM2[5539]<=26'd11156119; ROM3[5539]<=26'd9737634; ROM4[5539]<=26'd23443560;
ROM1[5540]<=26'd2008929; ROM2[5540]<=26'd11157229; ROM3[5540]<=26'd9732048; ROM4[5540]<=26'd23442957;
ROM1[5541]<=26'd2018455; ROM2[5541]<=26'd11162370; ROM3[5541]<=26'd9733049; ROM4[5541]<=26'd23446968;
ROM1[5542]<=26'd2016741; ROM2[5542]<=26'd11164344; ROM3[5542]<=26'd9739858; ROM4[5542]<=26'd23451131;
ROM1[5543]<=26'd2005604; ROM2[5543]<=26'd11160423; ROM3[5543]<=26'd9743616; ROM4[5543]<=26'd23450505;
ROM1[5544]<=26'd1995761; ROM2[5544]<=26'd11155693; ROM3[5544]<=26'd9743701; ROM4[5544]<=26'd23447168;
ROM1[5545]<=26'd1988047; ROM2[5545]<=26'd11151149; ROM3[5545]<=26'd9746128; ROM4[5545]<=26'd23446531;
ROM1[5546]<=26'd1985650; ROM2[5546]<=26'd11148651; ROM3[5546]<=26'd9746133; ROM4[5546]<=26'd23445085;
ROM1[5547]<=26'd1991752; ROM2[5547]<=26'd11150447; ROM3[5547]<=26'd9746167; ROM4[5547]<=26'd23446472;
ROM1[5548]<=26'd2005847; ROM2[5548]<=26'd11155683; ROM3[5548]<=26'd9744681; ROM4[5548]<=26'd23448692;
ROM1[5549]<=26'd2009620; ROM2[5549]<=26'd11153220; ROM3[5549]<=26'd9735365; ROM4[5549]<=26'd23444782;
ROM1[5550]<=26'd1997583; ROM2[5550]<=26'd11144965; ROM3[5550]<=26'd9729584; ROM4[5550]<=26'd23439680;
ROM1[5551]<=26'd1987833; ROM2[5551]<=26'd11140589; ROM3[5551]<=26'd9730901; ROM4[5551]<=26'd23436578;
ROM1[5552]<=26'd1979274; ROM2[5552]<=26'd11137189; ROM3[5552]<=26'd9731430; ROM4[5552]<=26'd23435240;
ROM1[5553]<=26'd1973269; ROM2[5553]<=26'd11138233; ROM3[5553]<=26'd9733947; ROM4[5553]<=26'd23436374;
ROM1[5554]<=26'd1974563; ROM2[5554]<=26'd11146695; ROM3[5554]<=26'd9742138; ROM4[5554]<=26'd23443688;
ROM1[5555]<=26'd1976715; ROM2[5555]<=26'd11148512; ROM3[5555]<=26'd9739665; ROM4[5555]<=26'd23444381;
ROM1[5556]<=26'd1985895; ROM2[5556]<=26'd11148586; ROM3[5556]<=26'd9733030; ROM4[5556]<=26'd23443681;
ROM1[5557]<=26'd2006228; ROM2[5557]<=26'd11154783; ROM3[5557]<=26'd9733973; ROM4[5557]<=26'd23450283;
ROM1[5558]<=26'd2016360; ROM2[5558]<=26'd11160875; ROM3[5558]<=26'd9739534; ROM4[5558]<=26'd23455375;
ROM1[5559]<=26'd2012114; ROM2[5559]<=26'd11161262; ROM3[5559]<=26'd9743194; ROM4[5559]<=26'd23457731;
ROM1[5560]<=26'd2006555; ROM2[5560]<=26'd11163017; ROM3[5560]<=26'd9749105; ROM4[5560]<=26'd23459720;
ROM1[5561]<=26'd2001081; ROM2[5561]<=26'd11163562; ROM3[5561]<=26'd9750401; ROM4[5561]<=26'd23456952;
ROM1[5562]<=26'd1990118; ROM2[5562]<=26'd11157417; ROM3[5562]<=26'd9743948; ROM4[5562]<=26'd23449589;
ROM1[5563]<=26'd1990909; ROM2[5563]<=26'd11157772; ROM3[5563]<=26'd9743545; ROM4[5563]<=26'd23448469;
ROM1[5564]<=26'd2001293; ROM2[5564]<=26'd11158975; ROM3[5564]<=26'd9740676; ROM4[5564]<=26'd23448818;
ROM1[5565]<=26'd2015494; ROM2[5565]<=26'd11162357; ROM3[5565]<=26'd9736536; ROM4[5565]<=26'd23451156;
ROM1[5566]<=26'd2023721; ROM2[5566]<=26'd11167305; ROM3[5566]<=26'd9739869; ROM4[5566]<=26'd23455293;
ROM1[5567]<=26'd2019092; ROM2[5567]<=26'd11166333; ROM3[5567]<=26'd9742415; ROM4[5567]<=26'd23455011;
ROM1[5568]<=26'd2011032; ROM2[5568]<=26'd11163360; ROM3[5568]<=26'd9744720; ROM4[5568]<=26'd23454400;
ROM1[5569]<=26'd2011226; ROM2[5569]<=26'd11167729; ROM3[5569]<=26'd9753879; ROM4[5569]<=26'd23460310;
ROM1[5570]<=26'd2014711; ROM2[5570]<=26'd11176452; ROM3[5570]<=26'd9764737; ROM4[5570]<=26'd23469707;
ROM1[5571]<=26'd2009672; ROM2[5571]<=26'd11173393; ROM3[5571]<=26'd9761468; ROM4[5571]<=26'd23467713;
ROM1[5572]<=26'd2010174; ROM2[5572]<=26'd11169059; ROM3[5572]<=26'd9755967; ROM4[5572]<=26'd23462951;
ROM1[5573]<=26'd2016363; ROM2[5573]<=26'd11163496; ROM3[5573]<=26'd9745927; ROM4[5573]<=26'd23457059;
ROM1[5574]<=26'd2021498; ROM2[5574]<=26'd11159199; ROM3[5574]<=26'd9739023; ROM4[5574]<=26'd23453254;
ROM1[5575]<=26'd2019186; ROM2[5575]<=26'd11158638; ROM3[5575]<=26'd9740993; ROM4[5575]<=26'd23454136;
ROM1[5576]<=26'd2012166; ROM2[5576]<=26'd11157236; ROM3[5576]<=26'd9745761; ROM4[5576]<=26'd23455203;
ROM1[5577]<=26'd2006986; ROM2[5577]<=26'd11156291; ROM3[5577]<=26'd9750176; ROM4[5577]<=26'd23455544;
ROM1[5578]<=26'd1999156; ROM2[5578]<=26'd11153205; ROM3[5578]<=26'd9749561; ROM4[5578]<=26'd23453338;
ROM1[5579]<=26'd1999361; ROM2[5579]<=26'd11156306; ROM3[5579]<=26'd9757233; ROM4[5579]<=26'd23457517;
ROM1[5580]<=26'd2008665; ROM2[5580]<=26'd11163643; ROM3[5580]<=26'd9763602; ROM4[5580]<=26'd23464821;
ROM1[5581]<=26'd2009769; ROM2[5581]<=26'd11158809; ROM3[5581]<=26'd9753784; ROM4[5581]<=26'd23457555;
ROM1[5582]<=26'd2009148; ROM2[5582]<=26'd11147745; ROM3[5582]<=26'd9739598; ROM4[5582]<=26'd23446192;
ROM1[5583]<=26'd2000413; ROM2[5583]<=26'd11139634; ROM3[5583]<=26'd9733272; ROM4[5583]<=26'd23438648;
ROM1[5584]<=26'd1987917; ROM2[5584]<=26'd11134796; ROM3[5584]<=26'd9732969; ROM4[5584]<=26'd23434257;
ROM1[5585]<=26'd1986295; ROM2[5585]<=26'd11137841; ROM3[5585]<=26'd9742209; ROM4[5585]<=26'd23440747;
ROM1[5586]<=26'd1981976; ROM2[5586]<=26'd11137052; ROM3[5586]<=26'd9745732; ROM4[5586]<=26'd23442210;
ROM1[5587]<=26'd1970587; ROM2[5587]<=26'd11130786; ROM3[5587]<=26'd9741704; ROM4[5587]<=26'd23435534;
ROM1[5588]<=26'd1968729; ROM2[5588]<=26'd11128064; ROM3[5588]<=26'd9740431; ROM4[5588]<=26'd23433577;
ROM1[5589]<=26'd1974760; ROM2[5589]<=26'd11126889; ROM3[5589]<=26'd9735008; ROM4[5589]<=26'd23432611;
ROM1[5590]<=26'd1986080; ROM2[5590]<=26'd11127262; ROM3[5590]<=26'd9728892; ROM4[5590]<=26'd23432937;
ROM1[5591]<=26'd1994440; ROM2[5591]<=26'd11130331; ROM3[5591]<=26'd9729809; ROM4[5591]<=26'd23438224;
ROM1[5592]<=26'd1994019; ROM2[5592]<=26'd11135806; ROM3[5592]<=26'd9735374; ROM4[5592]<=26'd23442756;
ROM1[5593]<=26'd1992520; ROM2[5593]<=26'd11142611; ROM3[5593]<=26'd9745473; ROM4[5593]<=26'd23448595;
ROM1[5594]<=26'd1982234; ROM2[5594]<=26'd11139604; ROM3[5594]<=26'd9745758; ROM4[5594]<=26'd23446340;
ROM1[5595]<=26'd1972366; ROM2[5595]<=26'd11136559; ROM3[5595]<=26'd9744149; ROM4[5595]<=26'd23443030;
ROM1[5596]<=26'd1970622; ROM2[5596]<=26'd11135418; ROM3[5596]<=26'd9740674; ROM4[5596]<=26'd23441485;
ROM1[5597]<=26'd1974927; ROM2[5597]<=26'd11133742; ROM3[5597]<=26'd9735354; ROM4[5597]<=26'd23440365;
ROM1[5598]<=26'd1994975; ROM2[5598]<=26'd11142137; ROM3[5598]<=26'd9738113; ROM4[5598]<=26'd23447491;
ROM1[5599]<=26'd2009884; ROM2[5599]<=26'd11148493; ROM3[5599]<=26'd9739427; ROM4[5599]<=26'd23452620;
ROM1[5600]<=26'd2008560; ROM2[5600]<=26'd11149690; ROM3[5600]<=26'd9743811; ROM4[5600]<=26'd23456535;
ROM1[5601]<=26'd2008207; ROM2[5601]<=26'd11156050; ROM3[5601]<=26'd9752826; ROM4[5601]<=26'd23463541;
ROM1[5602]<=26'd2007511; ROM2[5602]<=26'd11159351; ROM3[5602]<=26'd9757519; ROM4[5602]<=26'd23466395;
ROM1[5603]<=26'd1998549; ROM2[5603]<=26'd11156843; ROM3[5603]<=26'd9756291; ROM4[5603]<=26'd23463446;
ROM1[5604]<=26'd1991723; ROM2[5604]<=26'd11157350; ROM3[5604]<=26'd9755712; ROM4[5604]<=26'd23462488;
ROM1[5605]<=26'd1996186; ROM2[5605]<=26'd11159628; ROM3[5605]<=26'd9755392; ROM4[5605]<=26'd23463486;
ROM1[5606]<=26'd2004264; ROM2[5606]<=26'd11158074; ROM3[5606]<=26'd9749864; ROM4[5606]<=26'd23459483;
ROM1[5607]<=26'd2016426; ROM2[5607]<=26'd11160297; ROM3[5607]<=26'd9745679; ROM4[5607]<=26'd23461589;
ROM1[5608]<=26'd2018866; ROM2[5608]<=26'd11161308; ROM3[5608]<=26'd9746439; ROM4[5608]<=26'd23463594;
ROM1[5609]<=26'd2005939; ROM2[5609]<=26'd11154043; ROM3[5609]<=26'd9744151; ROM4[5609]<=26'd23457285;
ROM1[5610]<=26'd1999796; ROM2[5610]<=26'd11156318; ROM3[5610]<=26'd9749406; ROM4[5610]<=26'd23460554;
ROM1[5611]<=26'd2005308; ROM2[5611]<=26'd11168026; ROM3[5611]<=26'd9762588; ROM4[5611]<=26'd23471020;
ROM1[5612]<=26'd1998006; ROM2[5612]<=26'd11165558; ROM3[5612]<=26'd9761258; ROM4[5612]<=26'd23467315;
ROM1[5613]<=26'd1988713; ROM2[5613]<=26'd11156560; ROM3[5613]<=26'd9748850; ROM4[5613]<=26'd23455526;
ROM1[5614]<=26'd1999741; ROM2[5614]<=26'd11158770; ROM3[5614]<=26'd9746819; ROM4[5614]<=26'd23457256;
ROM1[5615]<=26'd2014649; ROM2[5615]<=26'd11159909; ROM3[5615]<=26'd9742230; ROM4[5615]<=26'd23458057;
ROM1[5616]<=26'd2012070; ROM2[5616]<=26'd11153047; ROM3[5616]<=26'd9733465; ROM4[5616]<=26'd23450250;
ROM1[5617]<=26'd2001649; ROM2[5617]<=26'd11150125; ROM3[5617]<=26'd9733493; ROM4[5617]<=26'd23448334;
ROM1[5618]<=26'd1988836; ROM2[5618]<=26'd11149119; ROM3[5618]<=26'd9733127; ROM4[5618]<=26'd23443987;
ROM1[5619]<=26'd1976126; ROM2[5619]<=26'd11143583; ROM3[5619]<=26'd9729040; ROM4[5619]<=26'd23436607;
ROM1[5620]<=26'd1971863; ROM2[5620]<=26'd11145295; ROM3[5620]<=26'd9730408; ROM4[5620]<=26'd23439570;
ROM1[5621]<=26'd1975861; ROM2[5621]<=26'd11149894; ROM3[5621]<=26'd9736143; ROM4[5621]<=26'd23443898;
ROM1[5622]<=26'd1981784; ROM2[5622]<=26'd11151360; ROM3[5622]<=26'd9736560; ROM4[5622]<=26'd23444982;
ROM1[5623]<=26'd1995373; ROM2[5623]<=26'd11154953; ROM3[5623]<=26'd9731721; ROM4[5623]<=26'd23446698;
ROM1[5624]<=26'd2005743; ROM2[5624]<=26'd11156922; ROM3[5624]<=26'd9728826; ROM4[5624]<=26'd23446634;
ROM1[5625]<=26'd1998146; ROM2[5625]<=26'd11152167; ROM3[5625]<=26'd9724921; ROM4[5625]<=26'd23443245;
ROM1[5626]<=26'd1989738; ROM2[5626]<=26'd11151247; ROM3[5626]<=26'd9726011; ROM4[5626]<=26'd23441947;
ROM1[5627]<=26'd1985121; ROM2[5627]<=26'd11152087; ROM3[5627]<=26'd9731962; ROM4[5627]<=26'd23443797;
ROM1[5628]<=26'd1978374; ROM2[5628]<=26'd11150683; ROM3[5628]<=26'd9735466; ROM4[5628]<=26'd23446789;
ROM1[5629]<=26'd1979003; ROM2[5629]<=26'd11155751; ROM3[5629]<=26'd9742907; ROM4[5629]<=26'd23453984;
ROM1[5630]<=26'd1986173; ROM2[5630]<=26'd11157325; ROM3[5630]<=26'd9745001; ROM4[5630]<=26'd23458747;
ROM1[5631]<=26'd1997545; ROM2[5631]<=26'd11156522; ROM3[5631]<=26'd9739720; ROM4[5631]<=26'd23458895;
ROM1[5632]<=26'd2009345; ROM2[5632]<=26'd11158644; ROM3[5632]<=26'd9736527; ROM4[5632]<=26'd23459534;
ROM1[5633]<=26'd2013429; ROM2[5633]<=26'd11163912; ROM3[5633]<=26'd9741260; ROM4[5633]<=26'd23464129;
ROM1[5634]<=26'd2014765; ROM2[5634]<=26'd11172441; ROM3[5634]<=26'd9752612; ROM4[5634]<=26'd23473259;
ROM1[5635]<=26'd2009691; ROM2[5635]<=26'd11172042; ROM3[5635]<=26'd9759324; ROM4[5635]<=26'd23476248;
ROM1[5636]<=26'd1999460; ROM2[5636]<=26'd11163655; ROM3[5636]<=26'd9755987; ROM4[5636]<=26'd23471003;
ROM1[5637]<=26'd1989110; ROM2[5637]<=26'd11155644; ROM3[5637]<=26'd9753393; ROM4[5637]<=26'd23466011;
ROM1[5638]<=26'd1982478; ROM2[5638]<=26'd11148339; ROM3[5638]<=26'd9747825; ROM4[5638]<=26'd23461240;
ROM1[5639]<=26'd1985160; ROM2[5639]<=26'd11145028; ROM3[5639]<=26'd9741102; ROM4[5639]<=26'd23456961;
ROM1[5640]<=26'd2002723; ROM2[5640]<=26'd11150181; ROM3[5640]<=26'd9741269; ROM4[5640]<=26'd23458768;
ROM1[5641]<=26'd2009473; ROM2[5641]<=26'd11153360; ROM3[5641]<=26'd9742458; ROM4[5641]<=26'd23463127;
ROM1[5642]<=26'd1995987; ROM2[5642]<=26'd11144810; ROM3[5642]<=26'd9739583; ROM4[5642]<=26'd23456616;
ROM1[5643]<=26'd1981352; ROM2[5643]<=26'd11136254; ROM3[5643]<=26'd9739076; ROM4[5643]<=26'd23450072;
ROM1[5644]<=26'd1975488; ROM2[5644]<=26'd11135413; ROM3[5644]<=26'd9741337; ROM4[5644]<=26'd23451411;
ROM1[5645]<=26'd1971452; ROM2[5645]<=26'd11135758; ROM3[5645]<=26'd9744640; ROM4[5645]<=26'd23452611;
ROM1[5646]<=26'd1970844; ROM2[5646]<=26'd11137963; ROM3[5646]<=26'd9746602; ROM4[5646]<=26'd23453259;
ROM1[5647]<=26'd1977382; ROM2[5647]<=26'd11141178; ROM3[5647]<=26'd9747032; ROM4[5647]<=26'd23455010;
ROM1[5648]<=26'd1987533; ROM2[5648]<=26'd11140660; ROM3[5648]<=26'd9743128; ROM4[5648]<=26'd23453443;
ROM1[5649]<=26'd1992616; ROM2[5649]<=26'd11136908; ROM3[5649]<=26'd9735935; ROM4[5649]<=26'd23449786;
ROM1[5650]<=26'd1993881; ROM2[5650]<=26'd11140828; ROM3[5650]<=26'd9739704; ROM4[5650]<=26'd23454555;
ROM1[5651]<=26'd1992384; ROM2[5651]<=26'd11146632; ROM3[5651]<=26'd9746774; ROM4[5651]<=26'd23461111;
ROM1[5652]<=26'd1982736; ROM2[5652]<=26'd11142867; ROM3[5652]<=26'd9747341; ROM4[5652]<=26'd23459360;
ROM1[5653]<=26'd1979744; ROM2[5653]<=26'd11145614; ROM3[5653]<=26'd9752423; ROM4[5653]<=26'd23461787;
ROM1[5654]<=26'd1979182; ROM2[5654]<=26'd11149033; ROM3[5654]<=26'd9755746; ROM4[5654]<=26'd23465002;
ROM1[5655]<=26'd1979025; ROM2[5655]<=26'd11148410; ROM3[5655]<=26'd9750843; ROM4[5655]<=26'd23460780;
ROM1[5656]<=26'd1990066; ROM2[5656]<=26'd11151878; ROM3[5656]<=26'd9745782; ROM4[5656]<=26'd23458274;
ROM1[5657]<=26'd2002824; ROM2[5657]<=26'd11154996; ROM3[5657]<=26'd9739345; ROM4[5657]<=26'd23457840;
ROM1[5658]<=26'd2000345; ROM2[5658]<=26'd11153615; ROM3[5658]<=26'd9734199; ROM4[5658]<=26'd23453659;
ROM1[5659]<=26'd1993134; ROM2[5659]<=26'd11153019; ROM3[5659]<=26'd9736392; ROM4[5659]<=26'd23453983;
ROM1[5660]<=26'd1987640; ROM2[5660]<=26'd11153918; ROM3[5660]<=26'd9741825; ROM4[5660]<=26'd23456454;
ROM1[5661]<=26'd1984629; ROM2[5661]<=26'd11157033; ROM3[5661]<=26'd9745390; ROM4[5661]<=26'd23458272;
ROM1[5662]<=26'd1984456; ROM2[5662]<=26'd11162754; ROM3[5662]<=26'd9752251; ROM4[5662]<=26'd23463726;
ROM1[5663]<=26'd1985433; ROM2[5663]<=26'd11162518; ROM3[5663]<=26'd9752212; ROM4[5663]<=26'd23463897;
ROM1[5664]<=26'd1993316; ROM2[5664]<=26'd11163102; ROM3[5664]<=26'd9747706; ROM4[5664]<=26'd23464970;
ROM1[5665]<=26'd2004798; ROM2[5665]<=26'd11164056; ROM3[5665]<=26'd9741800; ROM4[5665]<=26'd23464573;
ROM1[5666]<=26'd2003048; ROM2[5666]<=26'd11158304; ROM3[5666]<=26'd9734347; ROM4[5666]<=26'd23460889;
ROM1[5667]<=26'd1996734; ROM2[5667]<=26'd11156858; ROM3[5667]<=26'd9735106; ROM4[5667]<=26'd23461600;
ROM1[5668]<=26'd1990727; ROM2[5668]<=26'd11160466; ROM3[5668]<=26'd9740135; ROM4[5668]<=26'd23465245;
ROM1[5669]<=26'd1984877; ROM2[5669]<=26'd11160401; ROM3[5669]<=26'd9742373; ROM4[5669]<=26'd23465878;
ROM1[5670]<=26'd1977093; ROM2[5670]<=26'd11156308; ROM3[5670]<=26'd9742503; ROM4[5670]<=26'd23462648;
ROM1[5671]<=26'd1975986; ROM2[5671]<=26'd11155966; ROM3[5671]<=26'd9744060; ROM4[5671]<=26'd23463055;
ROM1[5672]<=26'd1987655; ROM2[5672]<=26'd11161720; ROM3[5672]<=26'd9747406; ROM4[5672]<=26'd23468347;
ROM1[5673]<=26'd2001521; ROM2[5673]<=26'd11164211; ROM3[5673]<=26'd9742927; ROM4[5673]<=26'd23467129;
ROM1[5674]<=26'd2008961; ROM2[5674]<=26'd11164144; ROM3[5674]<=26'd9736420; ROM4[5674]<=26'd23462656;
ROM1[5675]<=26'd2006713; ROM2[5675]<=26'd11164894; ROM3[5675]<=26'd9737626; ROM4[5675]<=26'd23462200;
ROM1[5676]<=26'd2001014; ROM2[5676]<=26'd11164772; ROM3[5676]<=26'd9742896; ROM4[5676]<=26'd23463459;
ROM1[5677]<=26'd2000226; ROM2[5677]<=26'd11167891; ROM3[5677]<=26'd9753575; ROM4[5677]<=26'd23469773;
ROM1[5678]<=26'd1993236; ROM2[5678]<=26'd11165347; ROM3[5678]<=26'd9756253; ROM4[5678]<=26'd23471050;
ROM1[5679]<=26'd1976469; ROM2[5679]<=26'd11151902; ROM3[5679]<=26'd9747614; ROM4[5679]<=26'd23460023;
ROM1[5680]<=26'd1976701; ROM2[5680]<=26'd11148045; ROM3[5680]<=26'd9742453; ROM4[5680]<=26'd23455568;
ROM1[5681]<=26'd1989907; ROM2[5681]<=26'd11153313; ROM3[5681]<=26'd9740290; ROM4[5681]<=26'd23457896;
ROM1[5682]<=26'd2005686; ROM2[5682]<=26'd11158499; ROM3[5682]<=26'd9740861; ROM4[5682]<=26'd23461149;
ROM1[5683]<=26'd2008127; ROM2[5683]<=26'd11160846; ROM3[5683]<=26'd9741987; ROM4[5683]<=26'd23463422;
ROM1[5684]<=26'd1994940; ROM2[5684]<=26'd11153595; ROM3[5684]<=26'd9740050; ROM4[5684]<=26'd23457475;
ROM1[5685]<=26'd1983891; ROM2[5685]<=26'd11146599; ROM3[5685]<=26'd9739742; ROM4[5685]<=26'd23454101;
ROM1[5686]<=26'd1985002; ROM2[5686]<=26'd11150901; ROM3[5686]<=26'd9747007; ROM4[5686]<=26'd23459778;
ROM1[5687]<=26'd1982556; ROM2[5687]<=26'd11154049; ROM3[5687]<=26'd9754302; ROM4[5687]<=26'd23463444;
ROM1[5688]<=26'd1977704; ROM2[5688]<=26'd11152529; ROM3[5688]<=26'd9751609; ROM4[5688]<=26'd23460018;
ROM1[5689]<=26'd1978762; ROM2[5689]<=26'd11149874; ROM3[5689]<=26'd9743738; ROM4[5689]<=26'd23454908;
ROM1[5690]<=26'd1981666; ROM2[5690]<=26'd11140584; ROM3[5690]<=26'd9729131; ROM4[5690]<=26'd23445996;
ROM1[5691]<=26'd1989632; ROM2[5691]<=26'd11144671; ROM3[5691]<=26'd9726827; ROM4[5691]<=26'd23447947;
ROM1[5692]<=26'd1992115; ROM2[5692]<=26'd11152494; ROM3[5692]<=26'd9734658; ROM4[5692]<=26'd23454718;
ROM1[5693]<=26'd1984272; ROM2[5693]<=26'd11150169; ROM3[5693]<=26'd9737264; ROM4[5693]<=26'd23454362;
ROM1[5694]<=26'd1977696; ROM2[5694]<=26'd11151897; ROM3[5694]<=26'd9741369; ROM4[5694]<=26'd23456100;
ROM1[5695]<=26'd1973251; ROM2[5695]<=26'd11153186; ROM3[5695]<=26'd9746632; ROM4[5695]<=26'd23459989;
ROM1[5696]<=26'd1974961; ROM2[5696]<=26'd11156606; ROM3[5696]<=26'd9749246; ROM4[5696]<=26'd23464114;
ROM1[5697]<=26'd1986006; ROM2[5697]<=26'd11161780; ROM3[5697]<=26'd9750238; ROM4[5697]<=26'd23466597;
ROM1[5698]<=26'd1999971; ROM2[5698]<=26'd11163709; ROM3[5698]<=26'd9746930; ROM4[5698]<=26'd23466783;
ROM1[5699]<=26'd2007048; ROM2[5699]<=26'd11165019; ROM3[5699]<=26'd9743138; ROM4[5699]<=26'd23467629;
ROM1[5700]<=26'd2000783; ROM2[5700]<=26'd11164252; ROM3[5700]<=26'd9742885; ROM4[5700]<=26'd23466834;
ROM1[5701]<=26'd1987968; ROM2[5701]<=26'd11159000; ROM3[5701]<=26'd9741768; ROM4[5701]<=26'd23463100;
ROM1[5702]<=26'd1984232; ROM2[5702]<=26'd11161253; ROM3[5702]<=26'd9747307; ROM4[5702]<=26'd23465541;
ROM1[5703]<=26'd1979039; ROM2[5703]<=26'd11161243; ROM3[5703]<=26'd9748413; ROM4[5703]<=26'd23462597;
ROM1[5704]<=26'd1968460; ROM2[5704]<=26'd11153023; ROM3[5704]<=26'd9743898; ROM4[5704]<=26'd23455368;
ROM1[5705]<=26'd1968944; ROM2[5705]<=26'd11151261; ROM3[5705]<=26'd9742179; ROM4[5705]<=26'd23454101;
ROM1[5706]<=26'd1977797; ROM2[5706]<=26'd11152764; ROM3[5706]<=26'd9735724; ROM4[5706]<=26'd23451861;
ROM1[5707]<=26'd1989871; ROM2[5707]<=26'd11155220; ROM3[5707]<=26'd9730744; ROM4[5707]<=26'd23451816;
ROM1[5708]<=26'd1989064; ROM2[5708]<=26'd11153434; ROM3[5708]<=26'd9726577; ROM4[5708]<=26'd23449516;
ROM1[5709]<=26'd1981363; ROM2[5709]<=26'd11152598; ROM3[5709]<=26'd9727305; ROM4[5709]<=26'd23449654;
ROM1[5710]<=26'd1977493; ROM2[5710]<=26'd11155089; ROM3[5710]<=26'd9735419; ROM4[5710]<=26'd23454299;
ROM1[5711]<=26'd1972263; ROM2[5711]<=26'd11154930; ROM3[5711]<=26'd9737545; ROM4[5711]<=26'd23453709;
ROM1[5712]<=26'd1968506; ROM2[5712]<=26'd11156290; ROM3[5712]<=26'd9740910; ROM4[5712]<=26'd23455623;
ROM1[5713]<=26'd1973390; ROM2[5713]<=26'd11162064; ROM3[5713]<=26'd9745505; ROM4[5713]<=26'd23460463;
ROM1[5714]<=26'd1980599; ROM2[5714]<=26'd11163913; ROM3[5714]<=26'd9742156; ROM4[5714]<=26'd23459123;
ROM1[5715]<=26'd1987714; ROM2[5715]<=26'd11159518; ROM3[5715]<=26'd9732896; ROM4[5715]<=26'd23454851;
ROM1[5716]<=26'd1989629; ROM2[5716]<=26'd11157551; ROM3[5716]<=26'd9727798; ROM4[5716]<=26'd23453221;
ROM1[5717]<=26'd1981800; ROM2[5717]<=26'd11155719; ROM3[5717]<=26'd9726792; ROM4[5717]<=26'd23451112;
ROM1[5718]<=26'd1971986; ROM2[5718]<=26'd11153843; ROM3[5718]<=26'd9726885; ROM4[5718]<=26'd23449115;
ROM1[5719]<=26'd1971925; ROM2[5719]<=26'd11157520; ROM3[5719]<=26'd9731888; ROM4[5719]<=26'd23454245;
ROM1[5720]<=26'd1971052; ROM2[5720]<=26'd11162708; ROM3[5720]<=26'd9740311; ROM4[5720]<=26'd23459648;
ROM1[5721]<=26'd1970870; ROM2[5721]<=26'd11164893; ROM3[5721]<=26'd9743669; ROM4[5721]<=26'd23461623;
ROM1[5722]<=26'd1972944; ROM2[5722]<=26'd11161062; ROM3[5722]<=26'd9738084; ROM4[5722]<=26'd23458043;
ROM1[5723]<=26'd1981491; ROM2[5723]<=26'd11158325; ROM3[5723]<=26'd9729792; ROM4[5723]<=26'd23453440;
ROM1[5724]<=26'd1988711; ROM2[5724]<=26'd11157304; ROM3[5724]<=26'd9722657; ROM4[5724]<=26'd23450795;
ROM1[5725]<=26'd1981067; ROM2[5725]<=26'd11152145; ROM3[5725]<=26'd9718708; ROM4[5725]<=26'd23447368;
ROM1[5726]<=26'd1975681; ROM2[5726]<=26'd11152234; ROM3[5726]<=26'd9724684; ROM4[5726]<=26'd23451437;
ROM1[5727]<=26'd1976804; ROM2[5727]<=26'd11157992; ROM3[5727]<=26'd9737042; ROM4[5727]<=26'd23458704;
ROM1[5728]<=26'd1970272; ROM2[5728]<=26'd11156199; ROM3[5728]<=26'd9740826; ROM4[5728]<=26'd23456919;
ROM1[5729]<=26'd1965928; ROM2[5729]<=26'd11153206; ROM3[5729]<=26'd9741119; ROM4[5729]<=26'd23454294;
ROM1[5730]<=26'd1971750; ROM2[5730]<=26'd11155167; ROM3[5730]<=26'd9742844; ROM4[5730]<=26'd23457164;
ROM1[5731]<=26'd1982010; ROM2[5731]<=26'd11156839; ROM3[5731]<=26'd9741785; ROM4[5731]<=26'd23459358;
ROM1[5732]<=26'd1989541; ROM2[5732]<=26'd11154834; ROM3[5732]<=26'd9737105; ROM4[5732]<=26'd23457134;
ROM1[5733]<=26'd1986463; ROM2[5733]<=26'd11150945; ROM3[5733]<=26'd9735060; ROM4[5733]<=26'd23455727;
ROM1[5734]<=26'd1980057; ROM2[5734]<=26'd11149552; ROM3[5734]<=26'd9736466; ROM4[5734]<=26'd23454992;
ROM1[5735]<=26'd1976694; ROM2[5735]<=26'd11153067; ROM3[5735]<=26'd9742561; ROM4[5735]<=26'd23458238;
ROM1[5736]<=26'd1979176; ROM2[5736]<=26'd11158436; ROM3[5736]<=26'd9751618; ROM4[5736]<=26'd23465808;
ROM1[5737]<=26'd1973877; ROM2[5737]<=26'd11158652; ROM3[5737]<=26'd9754608; ROM4[5737]<=26'd23465057;
ROM1[5738]<=26'd1968763; ROM2[5738]<=26'd11155059; ROM3[5738]<=26'd9749669; ROM4[5738]<=26'd23461059;
ROM1[5739]<=26'd1973613; ROM2[5739]<=26'd11151267; ROM3[5739]<=26'd9742751; ROM4[5739]<=26'd23457263;
ROM1[5740]<=26'd1986691; ROM2[5740]<=26'd11151983; ROM3[5740]<=26'd9737593; ROM4[5740]<=26'd23456899;
ROM1[5741]<=26'd1992649; ROM2[5741]<=26'd11157044; ROM3[5741]<=26'd9737423; ROM4[5741]<=26'd23459684;
ROM1[5742]<=26'd1989393; ROM2[5742]<=26'd11160411; ROM3[5742]<=26'd9740943; ROM4[5742]<=26'd23462076;
ROM1[5743]<=26'd1979469; ROM2[5743]<=26'd11158531; ROM3[5743]<=26'd9740674; ROM4[5743]<=26'd23459729;
ROM1[5744]<=26'd1971476; ROM2[5744]<=26'd11158276; ROM3[5744]<=26'd9741098; ROM4[5744]<=26'd23459620;
ROM1[5745]<=26'd1969091; ROM2[5745]<=26'd11157888; ROM3[5745]<=26'd9746194; ROM4[5745]<=26'd23462981;
ROM1[5746]<=26'd1967447; ROM2[5746]<=26'd11155105; ROM3[5746]<=26'd9746493; ROM4[5746]<=26'd23461141;
ROM1[5747]<=26'd1975231; ROM2[5747]<=26'd11159809; ROM3[5747]<=26'd9746996; ROM4[5747]<=26'd23464366;
ROM1[5748]<=26'd1985109; ROM2[5748]<=26'd11159097; ROM3[5748]<=26'd9740803; ROM4[5748]<=26'd23461423;
ROM1[5749]<=26'd1986377; ROM2[5749]<=26'd11152088; ROM3[5749]<=26'd9729875; ROM4[5749]<=26'd23454178;
ROM1[5750]<=26'd1987386; ROM2[5750]<=26'd11155259; ROM3[5750]<=26'd9736129; ROM4[5750]<=26'd23460115;
ROM1[5751]<=26'd1974218; ROM2[5751]<=26'd11147052; ROM3[5751]<=26'd9735544; ROM4[5751]<=26'd23456662;
ROM1[5752]<=26'd1959630; ROM2[5752]<=26'd11135878; ROM3[5752]<=26'd9730794; ROM4[5752]<=26'd23450095;
ROM1[5753]<=26'd1956812; ROM2[5753]<=26'd11138141; ROM3[5753]<=26'd9736739; ROM4[5753]<=26'd23453958;
ROM1[5754]<=26'd1954323; ROM2[5754]<=26'd11139640; ROM3[5754]<=26'd9739399; ROM4[5754]<=26'd23455917;
ROM1[5755]<=26'd1959932; ROM2[5755]<=26'd11140964; ROM3[5755]<=26'd9741392; ROM4[5755]<=26'd23457894;
ROM1[5756]<=26'd1972331; ROM2[5756]<=26'd11144810; ROM3[5756]<=26'd9740265; ROM4[5756]<=26'd23459471;
ROM1[5757]<=26'd1984589; ROM2[5757]<=26'd11146701; ROM3[5757]<=26'd9734887; ROM4[5757]<=26'd23460745;
ROM1[5758]<=26'd1983022; ROM2[5758]<=26'd11144090; ROM3[5758]<=26'd9731868; ROM4[5758]<=26'd23458047;
ROM1[5759]<=26'd1977257; ROM2[5759]<=26'd11143602; ROM3[5759]<=26'd9732604; ROM4[5759]<=26'd23456341;
ROM1[5760]<=26'd1973123; ROM2[5760]<=26'd11146257; ROM3[5760]<=26'd9737420; ROM4[5760]<=26'd23460931;
ROM1[5761]<=26'd1969229; ROM2[5761]<=26'd11147873; ROM3[5761]<=26'd9741481; ROM4[5761]<=26'd23461389;
ROM1[5762]<=26'd1963157; ROM2[5762]<=26'd11147905; ROM3[5762]<=26'd9742004; ROM4[5762]<=26'd23459061;
ROM1[5763]<=26'd1959752; ROM2[5763]<=26'd11145198; ROM3[5763]<=26'd9737268; ROM4[5763]<=26'd23455552;
ROM1[5764]<=26'd1965025; ROM2[5764]<=26'd11143907; ROM3[5764]<=26'd9732283; ROM4[5764]<=26'd23452011;
ROM1[5765]<=26'd1977420; ROM2[5765]<=26'd11147007; ROM3[5765]<=26'd9727744; ROM4[5765]<=26'd23451371;
ROM1[5766]<=26'd1978789; ROM2[5766]<=26'd11145859; ROM3[5766]<=26'd9723108; ROM4[5766]<=26'd23449952;
ROM1[5767]<=26'd1973717; ROM2[5767]<=26'd11145806; ROM3[5767]<=26'd9725405; ROM4[5767]<=26'd23450970;
ROM1[5768]<=26'd1969710; ROM2[5768]<=26'd11147110; ROM3[5768]<=26'd9728736; ROM4[5768]<=26'd23451621;
ROM1[5769]<=26'd1962694; ROM2[5769]<=26'd11143748; ROM3[5769]<=26'd9728405; ROM4[5769]<=26'd23448900;
ROM1[5770]<=26'd1957672; ROM2[5770]<=26'd11143990; ROM3[5770]<=26'd9731505; ROM4[5770]<=26'd23450092;
ROM1[5771]<=26'd1956655; ROM2[5771]<=26'd11145649; ROM3[5771]<=26'd9733790; ROM4[5771]<=26'd23452336;
ROM1[5772]<=26'd1971696; ROM2[5772]<=26'd11156964; ROM3[5772]<=26'd9741014; ROM4[5772]<=26'd23461923;
ROM1[5773]<=26'd1987628; ROM2[5773]<=26'd11162194; ROM3[5773]<=26'd9738647; ROM4[5773]<=26'd23465168;
ROM1[5774]<=26'd1987889; ROM2[5774]<=26'd11153980; ROM3[5774]<=26'd9727853; ROM4[5774]<=26'd23457781;
ROM1[5775]<=26'd1981773; ROM2[5775]<=26'd11151824; ROM3[5775]<=26'd9724983; ROM4[5775]<=26'd23454587;
ROM1[5776]<=26'd1975027; ROM2[5776]<=26'd11150915; ROM3[5776]<=26'd9728171; ROM4[5776]<=26'd23454999;
ROM1[5777]<=26'd1965538; ROM2[5777]<=26'd11144909; ROM3[5777]<=26'd9729259; ROM4[5777]<=26'd23451678;
ROM1[5778]<=26'd1960371; ROM2[5778]<=26'd11145627; ROM3[5778]<=26'd9730236; ROM4[5778]<=26'd23450741;
ROM1[5779]<=26'd1964535; ROM2[5779]<=26'd11152880; ROM3[5779]<=26'd9737732; ROM4[5779]<=26'd23458323;
ROM1[5780]<=26'd1963441; ROM2[5780]<=26'd11149220; ROM3[5780]<=26'd9733865; ROM4[5780]<=26'd23455824;
ROM1[5781]<=26'd1968665; ROM2[5781]<=26'd11143824; ROM3[5781]<=26'd9725216; ROM4[5781]<=26'd23450640;
ROM1[5782]<=26'd1984912; ROM2[5782]<=26'd11147020; ROM3[5782]<=26'd9725980; ROM4[5782]<=26'd23454970;
ROM1[5783]<=26'd1986133; ROM2[5783]<=26'd11149532; ROM3[5783]<=26'd9730100; ROM4[5783]<=26'd23457493;
ROM1[5784]<=26'd1982016; ROM2[5784]<=26'd11151596; ROM3[5784]<=26'd9734709; ROM4[5784]<=26'd23459996;
ROM1[5785]<=26'd1980350; ROM2[5785]<=26'd11155226; ROM3[5785]<=26'd9742463; ROM4[5785]<=26'd23464206;
ROM1[5786]<=26'd1975307; ROM2[5786]<=26'd11156303; ROM3[5786]<=26'd9747021; ROM4[5786]<=26'd23465952;
ROM1[5787]<=26'd1967505; ROM2[5787]<=26'd11154020; ROM3[5787]<=26'd9749318; ROM4[5787]<=26'd23464448;
ROM1[5788]<=26'd1971103; ROM2[5788]<=26'd11156653; ROM3[5788]<=26'd9755217; ROM4[5788]<=26'd23469885;
ROM1[5789]<=26'd1989362; ROM2[5789]<=26'd11166843; ROM3[5789]<=26'd9761436; ROM4[5789]<=26'd23481111;
ROM1[5790]<=26'd1998644; ROM2[5790]<=26'd11163387; ROM3[5790]<=26'd9751282; ROM4[5790]<=26'd23476512;
ROM1[5791]<=26'd1989850; ROM2[5791]<=26'd11149695; ROM3[5791]<=26'd9736378; ROM4[5791]<=26'd23462489;
ROM1[5792]<=26'd1983174; ROM2[5792]<=26'd11144983; ROM3[5792]<=26'd9735207; ROM4[5792]<=26'd23458782;
ROM1[5793]<=26'd1978369; ROM2[5793]<=26'd11146894; ROM3[5793]<=26'd9742638; ROM4[5793]<=26'd23463456;
ROM1[5794]<=26'd1979879; ROM2[5794]<=26'd11154353; ROM3[5794]<=26'd9753670; ROM4[5794]<=26'd23472679;
ROM1[5795]<=26'd1980271; ROM2[5795]<=26'd11159373; ROM3[5795]<=26'd9761820; ROM4[5795]<=26'd23479597;
ROM1[5796]<=26'd1977898; ROM2[5796]<=26'd11160519; ROM3[5796]<=26'd9761581; ROM4[5796]<=26'd23478094;
ROM1[5797]<=26'd1977528; ROM2[5797]<=26'd11156727; ROM3[5797]<=26'd9751387; ROM4[5797]<=26'd23470280;
ROM1[5798]<=26'd1987658; ROM2[5798]<=26'd11154763; ROM3[5798]<=26'd9743622; ROM4[5798]<=26'd23465589;
ROM1[5799]<=26'd1997445; ROM2[5799]<=26'd11156787; ROM3[5799]<=26'd9741351; ROM4[5799]<=26'd23467421;
ROM1[5800]<=26'd1992163; ROM2[5800]<=26'd11153227; ROM3[5800]<=26'd9740477; ROM4[5800]<=26'd23468462;
ROM1[5801]<=26'd1981128; ROM2[5801]<=26'd11147688; ROM3[5801]<=26'd9740540; ROM4[5801]<=26'd23464097;
ROM1[5802]<=26'd1975382; ROM2[5802]<=26'd11148669; ROM3[5802]<=26'd9743839; ROM4[5802]<=26'd23465662;
ROM1[5803]<=26'd1973721; ROM2[5803]<=26'd11151240; ROM3[5803]<=26'd9746610; ROM4[5803]<=26'd23468227;
ROM1[5804]<=26'd1966109; ROM2[5804]<=26'd11147795; ROM3[5804]<=26'd9745710; ROM4[5804]<=26'd23463884;
ROM1[5805]<=26'd1968054; ROM2[5805]<=26'd11146764; ROM3[5805]<=26'd9745138; ROM4[5805]<=26'd23464037;
ROM1[5806]<=26'd1975127; ROM2[5806]<=26'd11145173; ROM3[5806]<=26'd9739192; ROM4[5806]<=26'd23461038;
ROM1[5807]<=26'd1984671; ROM2[5807]<=26'd11146967; ROM3[5807]<=26'd9736012; ROM4[5807]<=26'd23462339;
ROM1[5808]<=26'd1983359; ROM2[5808]<=26'd11146552; ROM3[5808]<=26'd9736125; ROM4[5808]<=26'd23462266;
ROM1[5809]<=26'd1972724; ROM2[5809]<=26'd11142229; ROM3[5809]<=26'd9734140; ROM4[5809]<=26'd23459560;
ROM1[5810]<=26'd1965833; ROM2[5810]<=26'd11139933; ROM3[5810]<=26'd9735702; ROM4[5810]<=26'd23458475;
ROM1[5811]<=26'd1961583; ROM2[5811]<=26'd11138756; ROM3[5811]<=26'd9737436; ROM4[5811]<=26'd23457509;
ROM1[5812]<=26'd1956600; ROM2[5812]<=26'd11140671; ROM3[5812]<=26'd9737907; ROM4[5812]<=26'd23459541;
ROM1[5813]<=26'd1957048; ROM2[5813]<=26'd11142639; ROM3[5813]<=26'd9738854; ROM4[5813]<=26'd23459454;
ROM1[5814]<=26'd1966036; ROM2[5814]<=26'd11143268; ROM3[5814]<=26'd9736785; ROM4[5814]<=26'd23459375;
ROM1[5815]<=26'd1976589; ROM2[5815]<=26'd11141151; ROM3[5815]<=26'd9727868; ROM4[5815]<=26'd23456859;
ROM1[5816]<=26'd1981043; ROM2[5816]<=26'd11139827; ROM3[5816]<=26'd9724086; ROM4[5816]<=26'd23454035;
ROM1[5817]<=26'd1976505; ROM2[5817]<=26'd11141396; ROM3[5817]<=26'd9726382; ROM4[5817]<=26'd23454866;
ROM1[5818]<=26'd1969907; ROM2[5818]<=26'd11142713; ROM3[5818]<=26'd9731397; ROM4[5818]<=26'd23457844;
ROM1[5819]<=26'd1966318; ROM2[5819]<=26'd11144480; ROM3[5819]<=26'd9737224; ROM4[5819]<=26'd23460203;
ROM1[5820]<=26'd1954189; ROM2[5820]<=26'd11138298; ROM3[5820]<=26'd9732352; ROM4[5820]<=26'd23455026;
ROM1[5821]<=26'd1950370; ROM2[5821]<=26'd11135347; ROM3[5821]<=26'd9731304; ROM4[5821]<=26'd23453902;
ROM1[5822]<=26'd1957347; ROM2[5822]<=26'd11138047; ROM3[5822]<=26'd9730682; ROM4[5822]<=26'd23455438;
ROM1[5823]<=26'd1969782; ROM2[5823]<=26'd11139319; ROM3[5823]<=26'd9723653; ROM4[5823]<=26'd23453050;
ROM1[5824]<=26'd1981619; ROM2[5824]<=26'd11144545; ROM3[5824]<=26'd9725204; ROM4[5824]<=26'd23456093;
ROM1[5825]<=26'd1979705; ROM2[5825]<=26'd11149568; ROM3[5825]<=26'd9729898; ROM4[5825]<=26'd23458392;
ROM1[5826]<=26'd1973985; ROM2[5826]<=26'd11152101; ROM3[5826]<=26'd9736031; ROM4[5826]<=26'd23460755;
ROM1[5827]<=26'd1969801; ROM2[5827]<=26'd11152839; ROM3[5827]<=26'd9742138; ROM4[5827]<=26'd23463091;
ROM1[5828]<=26'd1968708; ROM2[5828]<=26'd11157368; ROM3[5828]<=26'd9748147; ROM4[5828]<=26'd23467040;
ROM1[5829]<=26'd1968054; ROM2[5829]<=26'd11157939; ROM3[5829]<=26'd9750086; ROM4[5829]<=26'd23468240;
ROM1[5830]<=26'd1969641; ROM2[5830]<=26'd11155444; ROM3[5830]<=26'd9747464; ROM4[5830]<=26'd23466875;
ROM1[5831]<=26'd1981116; ROM2[5831]<=26'd11159066; ROM3[5831]<=26'd9746040; ROM4[5831]<=26'd23467851;
ROM1[5832]<=26'd1995973; ROM2[5832]<=26'd11162383; ROM3[5832]<=26'd9743489; ROM4[5832]<=26'd23469486;
ROM1[5833]<=26'd1992084; ROM2[5833]<=26'd11158021; ROM3[5833]<=26'd9738264; ROM4[5833]<=26'd23465739;
ROM1[5834]<=26'd1981854; ROM2[5834]<=26'd11154582; ROM3[5834]<=26'd9738028; ROM4[5834]<=26'd23463778;
ROM1[5835]<=26'd1975178; ROM2[5835]<=26'd11154764; ROM3[5835]<=26'd9742900; ROM4[5835]<=26'd23466004;
ROM1[5836]<=26'd1969384; ROM2[5836]<=26'd11154025; ROM3[5836]<=26'd9744549; ROM4[5836]<=26'd23466288;
ROM1[5837]<=26'd1966778; ROM2[5837]<=26'd11154456; ROM3[5837]<=26'd9748217; ROM4[5837]<=26'd23467154;
ROM1[5838]<=26'd1969446; ROM2[5838]<=26'd11156852; ROM3[5838]<=26'd9748128; ROM4[5838]<=26'd23466829;
ROM1[5839]<=26'd1972545; ROM2[5839]<=26'd11151882; ROM3[5839]<=26'd9737838; ROM4[5839]<=26'd23461428;
ROM1[5840]<=26'd1984079; ROM2[5840]<=26'd11150350; ROM3[5840]<=26'd9732795; ROM4[5840]<=26'd23459221;
ROM1[5841]<=26'd1998660; ROM2[5841]<=26'd11163039; ROM3[5841]<=26'd9742175; ROM4[5841]<=26'd23470216;
ROM1[5842]<=26'd1996474; ROM2[5842]<=26'd11166554; ROM3[5842]<=26'd9747055; ROM4[5842]<=26'd23474517;
ROM1[5843]<=26'd1983178; ROM2[5843]<=26'd11161518; ROM3[5843]<=26'd9746319; ROM4[5843]<=26'd23470037;
ROM1[5844]<=26'd1970182; ROM2[5844]<=26'd11154093; ROM3[5844]<=26'd9742946; ROM4[5844]<=26'd23461999;
ROM1[5845]<=26'd1952788; ROM2[5845]<=26'd11141118; ROM3[5845]<=26'd9735910; ROM4[5845]<=26'd23450443;
ROM1[5846]<=26'd1949130; ROM2[5846]<=26'd11138065; ROM3[5846]<=26'd9735276; ROM4[5846]<=26'd23447618;
ROM1[5847]<=26'd1961432; ROM2[5847]<=26'd11144129; ROM3[5847]<=26'd9738899; ROM4[5847]<=26'd23452366;
ROM1[5848]<=26'd1977198; ROM2[5848]<=26'd11149405; ROM3[5848]<=26'd9737468; ROM4[5848]<=26'd23455021;
ROM1[5849]<=26'd1986783; ROM2[5849]<=26'd11151244; ROM3[5849]<=26'd9732958; ROM4[5849]<=26'd23455717;
ROM1[5850]<=26'd1983423; ROM2[5850]<=26'd11151870; ROM3[5850]<=26'd9732045; ROM4[5850]<=26'd23455432;
ROM1[5851]<=26'd1975650; ROM2[5851]<=26'd11150647; ROM3[5851]<=26'd9734137; ROM4[5851]<=26'd23453114;
ROM1[5852]<=26'd1969786; ROM2[5852]<=26'd11147072; ROM3[5852]<=26'd9736744; ROM4[5852]<=26'd23452199;
ROM1[5853]<=26'd1964219; ROM2[5853]<=26'd11145383; ROM3[5853]<=26'd9740739; ROM4[5853]<=26'd23454933;
ROM1[5854]<=26'd1957663; ROM2[5854]<=26'd11143658; ROM3[5854]<=26'd9740952; ROM4[5854]<=26'd23454020;
ROM1[5855]<=26'd1959987; ROM2[5855]<=26'd11145606; ROM3[5855]<=26'd9737376; ROM4[5855]<=26'd23453481;
ROM1[5856]<=26'd1975260; ROM2[5856]<=26'd11151666; ROM3[5856]<=26'd9734153; ROM4[5856]<=26'd23455066;
ROM1[5857]<=26'd1988473; ROM2[5857]<=26'd11154917; ROM3[5857]<=26'd9727875; ROM4[5857]<=26'd23454432;
ROM1[5858]<=26'd1983930; ROM2[5858]<=26'd11151890; ROM3[5858]<=26'd9724332; ROM4[5858]<=26'd23451274;
ROM1[5859]<=26'd1975419; ROM2[5859]<=26'd11149772; ROM3[5859]<=26'd9726008; ROM4[5859]<=26'd23449850;
ROM1[5860]<=26'd1970188; ROM2[5860]<=26'd11149139; ROM3[5860]<=26'd9729234; ROM4[5860]<=26'd23451853;
ROM1[5861]<=26'd1971453; ROM2[5861]<=26'd11150945; ROM3[5861]<=26'd9733369; ROM4[5861]<=26'd23454302;
ROM1[5862]<=26'd1970404; ROM2[5862]<=26'd11150751; ROM3[5862]<=26'd9737665; ROM4[5862]<=26'd23455571;
ROM1[5863]<=26'd1975887; ROM2[5863]<=26'd11152083; ROM3[5863]<=26'd9743234; ROM4[5863]<=26'd23460664;
ROM1[5864]<=26'd1990065; ROM2[5864]<=26'd11160400; ROM3[5864]<=26'd9746658; ROM4[5864]<=26'd23467645;
ROM1[5865]<=26'd1999854; ROM2[5865]<=26'd11160758; ROM3[5865]<=26'd9738901; ROM4[5865]<=26'd23465557;
ROM1[5866]<=26'd2003889; ROM2[5866]<=26'd11158589; ROM3[5866]<=26'd9733950; ROM4[5866]<=26'd23462440;
ROM1[5867]<=26'd2002385; ROM2[5867]<=26'd11161901; ROM3[5867]<=26'd9736485; ROM4[5867]<=26'd23463725;
ROM1[5868]<=26'd1990154; ROM2[5868]<=26'd11159954; ROM3[5868]<=26'd9738590; ROM4[5868]<=26'd23462470;
ROM1[5869]<=26'd1991980; ROM2[5869]<=26'd11164584; ROM3[5869]<=26'd9748257; ROM4[5869]<=26'd23468061;
ROM1[5870]<=26'd1998750; ROM2[5870]<=26'd11171074; ROM3[5870]<=26'd9754971; ROM4[5870]<=26'd23474341;
ROM1[5871]<=26'd1998989; ROM2[5871]<=26'd11165200; ROM3[5871]<=26'd9749046; ROM4[5871]<=26'd23468957;
ROM1[5872]<=26'd2008834; ROM2[5872]<=26'd11162679; ROM3[5872]<=26'd9741184; ROM4[5872]<=26'd23465443;
ROM1[5873]<=26'd2025151; ROM2[5873]<=26'd11166464; ROM3[5873]<=26'd9734833; ROM4[5873]<=26'd23466026;
ROM1[5874]<=26'd2045556; ROM2[5874]<=26'd11176836; ROM3[5874]<=26'd9739109; ROM4[5874]<=26'd23474382;
ROM1[5875]<=26'd2055829; ROM2[5875]<=26'd11186731; ROM3[5875]<=26'd9750046; ROM4[5875]<=26'd23485932;
ROM1[5876]<=26'd2052435; ROM2[5876]<=26'd11184340; ROM3[5876]<=26'd9752899; ROM4[5876]<=26'd23487961;
ROM1[5877]<=26'd2048893; ROM2[5877]<=26'd11180247; ROM3[5877]<=26'd9751917; ROM4[5877]<=26'd23485331;
ROM1[5878]<=26'd2048637; ROM2[5878]<=26'd11179777; ROM3[5878]<=26'd9753443; ROM4[5878]<=26'd23485507;
ROM1[5879]<=26'd2053138; ROM2[5879]<=26'd11182158; ROM3[5879]<=26'd9756443; ROM4[5879]<=26'd23488160;
ROM1[5880]<=26'd2070255; ROM2[5880]<=26'd11192959; ROM3[5880]<=26'd9763727; ROM4[5880]<=26'd23496403;
ROM1[5881]<=26'd2084389; ROM2[5881]<=26'd11195192; ROM3[5881]<=26'd9760599; ROM4[5881]<=26'd23497053;
ROM1[5882]<=26'd2091698; ROM2[5882]<=26'd11188833; ROM3[5882]<=26'd9748148; ROM4[5882]<=26'd23489779;
ROM1[5883]<=26'd2095907; ROM2[5883]<=26'd11189648; ROM3[5883]<=26'd9748551; ROM4[5883]<=26'd23490669;
ROM1[5884]<=26'd2094725; ROM2[5884]<=26'd11190016; ROM3[5884]<=26'd9752141; ROM4[5884]<=26'd23490970;
ROM1[5885]<=26'd2092074; ROM2[5885]<=26'd11189239; ROM3[5885]<=26'd9756263; ROM4[5885]<=26'd23491451;
ROM1[5886]<=26'd2092282; ROM2[5886]<=26'd11191319; ROM3[5886]<=26'd9760847; ROM4[5886]<=26'd23494120;
ROM1[5887]<=26'd2090525; ROM2[5887]<=26'd11191346; ROM3[5887]<=26'd9761229; ROM4[5887]<=26'd23494269;
ROM1[5888]<=26'd2095646; ROM2[5888]<=26'd11193299; ROM3[5888]<=26'd9759601; ROM4[5888]<=26'd23496536;
ROM1[5889]<=26'd2111867; ROM2[5889]<=26'd11200089; ROM3[5889]<=26'd9760156; ROM4[5889]<=26'd23501033;
ROM1[5890]<=26'd2129834; ROM2[5890]<=26'd11206147; ROM3[5890]<=26'd9758589; ROM4[5890]<=26'd23503770;
ROM1[5891]<=26'd2136980; ROM2[5891]<=26'd11210664; ROM3[5891]<=26'd9759824; ROM4[5891]<=26'd23506882;
ROM1[5892]<=26'd2134553; ROM2[5892]<=26'd11212815; ROM3[5892]<=26'd9764374; ROM4[5892]<=26'd23510064;
ROM1[5893]<=26'd2127003; ROM2[5893]<=26'd11210688; ROM3[5893]<=26'd9766751; ROM4[5893]<=26'd23509254;
ROM1[5894]<=26'd2116507; ROM2[5894]<=26'd11205019; ROM3[5894]<=26'd9763834; ROM4[5894]<=26'd23503992;
ROM1[5895]<=26'd2106974; ROM2[5895]<=26'd11200152; ROM3[5895]<=26'd9760239; ROM4[5895]<=26'd23497968;
ROM1[5896]<=26'd2106389; ROM2[5896]<=26'd11199964; ROM3[5896]<=26'd9760341; ROM4[5896]<=26'd23497639;
ROM1[5897]<=26'd2118707; ROM2[5897]<=26'd11205865; ROM3[5897]<=26'd9762693; ROM4[5897]<=26'd23503376;
ROM1[5898]<=26'd2135208; ROM2[5898]<=26'd11210698; ROM3[5898]<=26'd9764934; ROM4[5898]<=26'd23508450;
ROM1[5899]<=26'd2142165; ROM2[5899]<=26'd11210829; ROM3[5899]<=26'd9763671; ROM4[5899]<=26'd23509053;
ROM1[5900]<=26'd2133662; ROM2[5900]<=26'd11206660; ROM3[5900]<=26'd9761872; ROM4[5900]<=26'd23504500;
ROM1[5901]<=26'd2118552; ROM2[5901]<=26'd11200841; ROM3[5901]<=26'd9760238; ROM4[5901]<=26'd23499366;
ROM1[5902]<=26'd2108513; ROM2[5902]<=26'd11198785; ROM3[5902]<=26'd9761237; ROM4[5902]<=26'd23498297;
ROM1[5903]<=26'd2103008; ROM2[5903]<=26'd11197431; ROM3[5903]<=26'd9764308; ROM4[5903]<=26'd23499131;
ROM1[5904]<=26'd2094893; ROM2[5904]<=26'd11195044; ROM3[5904]<=26'd9764666; ROM4[5904]<=26'd23496665;
ROM1[5905]<=26'd2092780; ROM2[5905]<=26'd11193861; ROM3[5905]<=26'd9761439; ROM4[5905]<=26'd23493584;
ROM1[5906]<=26'd2103368; ROM2[5906]<=26'd11196810; ROM3[5906]<=26'd9758293; ROM4[5906]<=26'd23494595;
ROM1[5907]<=26'd2112527; ROM2[5907]<=26'd11198199; ROM3[5907]<=26'd9752107; ROM4[5907]<=26'd23493640;
ROM1[5908]<=26'd2109361; ROM2[5908]<=26'd11197126; ROM3[5908]<=26'd9750079; ROM4[5908]<=26'd23493472;
ROM1[5909]<=26'd2098189; ROM2[5909]<=26'd11194230; ROM3[5909]<=26'd9751636; ROM4[5909]<=26'd23492045;
ROM1[5910]<=26'd2089538; ROM2[5910]<=26'd11192152; ROM3[5910]<=26'd9753391; ROM4[5910]<=26'd23489437;
ROM1[5911]<=26'd2090155; ROM2[5911]<=26'd11199861; ROM3[5911]<=26'd9762725; ROM4[5911]<=26'd23497825;
ROM1[5912]<=26'd2090793; ROM2[5912]<=26'd11208532; ROM3[5912]<=26'd9772950; ROM4[5912]<=26'd23506285;
ROM1[5913]<=26'd2072362; ROM2[5913]<=26'd11192608; ROM3[5913]<=26'd9757331; ROM4[5913]<=26'd23490677;
ROM1[5914]<=26'd2061907; ROM2[5914]<=26'd11179572; ROM3[5914]<=26'd9740130; ROM4[5914]<=26'd23478643;
ROM1[5915]<=26'd2076387; ROM2[5915]<=26'd11183831; ROM3[5915]<=26'd9737167; ROM4[5915]<=26'd23480399;
ROM1[5916]<=26'd2078331; ROM2[5916]<=26'd11180708; ROM3[5916]<=26'd9733197; ROM4[5916]<=26'd23477501;
ROM1[5917]<=26'd2081159; ROM2[5917]<=26'd11188175; ROM3[5917]<=26'd9744877; ROM4[5917]<=26'd23486608;
ROM1[5918]<=26'd2078218; ROM2[5918]<=26'd11193390; ROM3[5918]<=26'd9755617; ROM4[5918]<=26'd23494830;
ROM1[5919]<=26'd2056379; ROM2[5919]<=26'd11179705; ROM3[5919]<=26'd9747092; ROM4[5919]<=26'd23482526;
ROM1[5920]<=26'd2042906; ROM2[5920]<=26'd11174488; ROM3[5920]<=26'd9744653; ROM4[5920]<=26'd23476786;
ROM1[5921]<=26'd2051575; ROM2[5921]<=26'd11183237; ROM3[5921]<=26'd9755542; ROM4[5921]<=26'd23487160;
ROM1[5922]<=26'd2056566; ROM2[5922]<=26'd11182960; ROM3[5922]<=26'd9753411; ROM4[5922]<=26'd23485695;
ROM1[5923]<=26'd2058474; ROM2[5923]<=26'd11177865; ROM3[5923]<=26'd9742336; ROM4[5923]<=26'd23478179;
ROM1[5924]<=26'd2060377; ROM2[5924]<=26'd11173458; ROM3[5924]<=26'd9737930; ROM4[5924]<=26'd23476259;
ROM1[5925]<=26'd2053590; ROM2[5925]<=26'd11170488; ROM3[5925]<=26'd9738153; ROM4[5925]<=26'd23475319;
ROM1[5926]<=26'd2051101; ROM2[5926]<=26'd11176609; ROM3[5926]<=26'd9747526; ROM4[5926]<=26'd23482597;
ROM1[5927]<=26'd2047249; ROM2[5927]<=26'd11178195; ROM3[5927]<=26'd9756435; ROM4[5927]<=26'd23486778;
ROM1[5928]<=26'd2036887; ROM2[5928]<=26'd11173320; ROM3[5928]<=26'd9757273; ROM4[5928]<=26'd23483112;
ROM1[5929]<=26'd2029138; ROM2[5929]<=26'd11171679; ROM3[5929]<=26'd9756779; ROM4[5929]<=26'd23481541;
ROM1[5930]<=26'd2033805; ROM2[5930]<=26'd11172753; ROM3[5930]<=26'd9761159; ROM4[5930]<=26'd23484179;
ROM1[5931]<=26'd2049193; ROM2[5931]<=26'd11178847; ROM3[5931]<=26'd9763395; ROM4[5931]<=26'd23490992;
ROM1[5932]<=26'd2052786; ROM2[5932]<=26'd11175128; ROM3[5932]<=26'd9752555; ROM4[5932]<=26'd23485717;
ROM1[5933]<=26'd2045867; ROM2[5933]<=26'd11169543; ROM3[5933]<=26'd9747685; ROM4[5933]<=26'd23479905;
ROM1[5934]<=26'd2036613; ROM2[5934]<=26'd11168068; ROM3[5934]<=26'd9748401; ROM4[5934]<=26'd23477584;
ROM1[5935]<=26'd2026020; ROM2[5935]<=26'd11164685; ROM3[5935]<=26'd9748849; ROM4[5935]<=26'd23475079;
ROM1[5936]<=26'd2023609; ROM2[5936]<=26'd11167879; ROM3[5936]<=26'd9755437; ROM4[5936]<=26'd23480204;
ROM1[5937]<=26'd2016878; ROM2[5937]<=26'd11166737; ROM3[5937]<=26'd9757953; ROM4[5937]<=26'd23480744;
ROM1[5938]<=26'd2009345; ROM2[5938]<=26'd11160410; ROM3[5938]<=26'd9750759; ROM4[5938]<=26'd23473456;
ROM1[5939]<=26'd2010735; ROM2[5939]<=26'd11154810; ROM3[5939]<=26'd9742579; ROM4[5939]<=26'd23469099;
ROM1[5940]<=26'd2025970; ROM2[5940]<=26'd11157766; ROM3[5940]<=26'd9739956; ROM4[5940]<=26'd23471720;
ROM1[5941]<=26'd2033629; ROM2[5941]<=26'd11161242; ROM3[5941]<=26'd9742309; ROM4[5941]<=26'd23475373;
ROM1[5942]<=26'd2033723; ROM2[5942]<=26'd11164751; ROM3[5942]<=26'd9747939; ROM4[5942]<=26'd23480703;
ROM1[5943]<=26'd2020579; ROM2[5943]<=26'd11157643; ROM3[5943]<=26'd9744902; ROM4[5943]<=26'd23473847;
ROM1[5944]<=26'd2005704; ROM2[5944]<=26'd11147810; ROM3[5944]<=26'd9739581; ROM4[5944]<=26'd23465611;
ROM1[5945]<=26'd1998999; ROM2[5945]<=26'd11147029; ROM3[5945]<=26'd9741207; ROM4[5945]<=26'd23466029;
ROM1[5946]<=26'd1991950; ROM2[5946]<=26'd11143200; ROM3[5946]<=26'd9740362; ROM4[5946]<=26'd23461584;
ROM1[5947]<=26'd1997823; ROM2[5947]<=26'd11143976; ROM3[5947]<=26'd9740638; ROM4[5947]<=26'd23462104;
ROM1[5948]<=26'd2014003; ROM2[5948]<=26'd11149174; ROM3[5948]<=26'd9739053; ROM4[5948]<=26'd23466499;
ROM1[5949]<=26'd2016868; ROM2[5949]<=26'd11148005; ROM3[5949]<=26'd9731311; ROM4[5949]<=26'd23462267;
ROM1[5950]<=26'd2009325; ROM2[5950]<=26'd11144742; ROM3[5950]<=26'd9727653; ROM4[5950]<=26'd23459299;
ROM1[5951]<=26'd2005492; ROM2[5951]<=26'd11147991; ROM3[5951]<=26'd9734161; ROM4[5951]<=26'd23463968;
ROM1[5952]<=26'd2004342; ROM2[5952]<=26'd11155458; ROM3[5952]<=26'd9744922; ROM4[5952]<=26'd23471663;
ROM1[5953]<=26'd1998045; ROM2[5953]<=26'd11156272; ROM3[5953]<=26'd9746957; ROM4[5953]<=26'd23471223;
ROM1[5954]<=26'd1987415; ROM2[5954]<=26'd11149635; ROM3[5954]<=26'd9741225; ROM4[5954]<=26'd23464139;
ROM1[5955]<=26'd1987174; ROM2[5955]<=26'd11148141; ROM3[5955]<=26'd9737835; ROM4[5955]<=26'd23461480;
ROM1[5956]<=26'd1995634; ROM2[5956]<=26'd11147144; ROM3[5956]<=26'd9731959; ROM4[5956]<=26'd23457592;
ROM1[5957]<=26'd2008472; ROM2[5957]<=26'd11148920; ROM3[5957]<=26'd9728312; ROM4[5957]<=26'd23457678;
ROM1[5958]<=26'd2011329; ROM2[5958]<=26'd11150950; ROM3[5958]<=26'd9729839; ROM4[5958]<=26'd23460136;
ROM1[5959]<=26'd2002387; ROM2[5959]<=26'd11151121; ROM3[5959]<=26'd9727745; ROM4[5959]<=26'd23458464;
ROM1[5960]<=26'd1992834; ROM2[5960]<=26'd11149736; ROM3[5960]<=26'd9727694; ROM4[5960]<=26'd23455056;
ROM1[5961]<=26'd1986360; ROM2[5961]<=26'd11147824; ROM3[5961]<=26'd9730320; ROM4[5961]<=26'd23454582;
ROM1[5962]<=26'd1982536; ROM2[5962]<=26'd11148984; ROM3[5962]<=26'd9734087; ROM4[5962]<=26'd23456627;
ROM1[5963]<=26'd1987619; ROM2[5963]<=26'd11152422; ROM3[5963]<=26'd9738422; ROM4[5963]<=26'd23459820;
ROM1[5964]<=26'd1997934; ROM2[5964]<=26'd11155220; ROM3[5964]<=26'd9736066; ROM4[5964]<=26'd23460656;
ROM1[5965]<=26'd2005288; ROM2[5965]<=26'd11151090; ROM3[5965]<=26'd9724894; ROM4[5965]<=26'd23454846;
ROM1[5966]<=26'd2005687; ROM2[5966]<=26'd11148394; ROM3[5966]<=26'd9721686; ROM4[5966]<=26'd23451979;
ROM1[5967]<=26'd1997296; ROM2[5967]<=26'd11145087; ROM3[5967]<=26'd9722239; ROM4[5967]<=26'd23449445;
ROM1[5968]<=26'd1987009; ROM2[5968]<=26'd11140953; ROM3[5968]<=26'd9722647; ROM4[5968]<=26'd23447886;
ROM1[5969]<=26'd1983393; ROM2[5969]<=26'd11142454; ROM3[5969]<=26'd9728675; ROM4[5969]<=26'd23451357;
ROM1[5970]<=26'd1980793; ROM2[5970]<=26'd11145394; ROM3[5970]<=26'd9738707; ROM4[5970]<=26'd23457627;
ROM1[5971]<=26'd1980350; ROM2[5971]<=26'd11143872; ROM3[5971]<=26'd9738479; ROM4[5971]<=26'd23457846;
ROM1[5972]<=26'd1982627; ROM2[5972]<=26'd11139883; ROM3[5972]<=26'd9733045; ROM4[5972]<=26'd23454082;
ROM1[5973]<=26'd1992845; ROM2[5973]<=26'd11140336; ROM3[5973]<=26'd9727825; ROM4[5973]<=26'd23453112;
ROM1[5974]<=26'd1999473; ROM2[5974]<=26'd11139953; ROM3[5974]<=26'd9721575; ROM4[5974]<=26'd23450925;
ROM1[5975]<=26'd1993143; ROM2[5975]<=26'd11138443; ROM3[5975]<=26'd9723293; ROM4[5975]<=26'd23450070;
ROM1[5976]<=26'd1985796; ROM2[5976]<=26'd11137212; ROM3[5976]<=26'd9726174; ROM4[5976]<=26'd23448536;
ROM1[5977]<=26'd1982997; ROM2[5977]<=26'd11138726; ROM3[5977]<=26'd9730295; ROM4[5977]<=26'd23448760;
ROM1[5978]<=26'd1979197; ROM2[5978]<=26'd11140642; ROM3[5978]<=26'd9734380; ROM4[5978]<=26'd23453157;
ROM1[5979]<=26'd1975454; ROM2[5979]<=26'd11140720; ROM3[5979]<=26'd9735803; ROM4[5979]<=26'd23453662;
ROM1[5980]<=26'd1981535; ROM2[5980]<=26'd11145337; ROM3[5980]<=26'd9736998; ROM4[5980]<=26'd23455499;
ROM1[5981]<=26'd2008222; ROM2[5981]<=26'd11161187; ROM3[5981]<=26'd9747294; ROM4[5981]<=26'd23470790;
ROM1[5982]<=26'd2021400; ROM2[5982]<=26'd11164350; ROM3[5982]<=26'd9742781; ROM4[5982]<=26'd23470301;
ROM1[5983]<=26'd2005982; ROM2[5983]<=26'd11148975; ROM3[5983]<=26'd9728040; ROM4[5983]<=26'd23456462;
ROM1[5984]<=26'd1996128; ROM2[5984]<=26'd11145788; ROM3[5984]<=26'd9729521; ROM4[5984]<=26'd23454701;
ROM1[5985]<=26'd1986491; ROM2[5985]<=26'd11145182; ROM3[5985]<=26'd9731550; ROM4[5985]<=26'd23453254;
ROM1[5986]<=26'd1977313; ROM2[5986]<=26'd11140510; ROM3[5986]<=26'd9729732; ROM4[5986]<=26'd23450099;
ROM1[5987]<=26'd1975554; ROM2[5987]<=26'd11142420; ROM3[5987]<=26'd9734979; ROM4[5987]<=26'd23452860;
ROM1[5988]<=26'd1979998; ROM2[5988]<=26'd11143913; ROM3[5988]<=26'd9738892; ROM4[5988]<=26'd23458005;
ROM1[5989]<=26'd1984189; ROM2[5989]<=26'd11139658; ROM3[5989]<=26'd9731864; ROM4[5989]<=26'd23454754;
ROM1[5990]<=26'd1996125; ROM2[5990]<=26'd11138593; ROM3[5990]<=26'd9724498; ROM4[5990]<=26'd23454157;
ROM1[5991]<=26'd2003642; ROM2[5991]<=26'd11142912; ROM3[5991]<=26'd9725553; ROM4[5991]<=26'd23459501;
ROM1[5992]<=26'd2004511; ROM2[5992]<=26'd11149936; ROM3[5992]<=26'd9734356; ROM4[5992]<=26'd23466046;
ROM1[5993]<=26'd1989730; ROM2[5993]<=26'd11141818; ROM3[5993]<=26'd9730543; ROM4[5993]<=26'd23460842;
ROM1[5994]<=26'd1973141; ROM2[5994]<=26'd11131546; ROM3[5994]<=26'd9722684; ROM4[5994]<=26'd23451383;
ROM1[5995]<=26'd1972712; ROM2[5995]<=26'd11137343; ROM3[5995]<=26'd9732126; ROM4[5995]<=26'd23457509;
ROM1[5996]<=26'd1971311; ROM2[5996]<=26'd11138267; ROM3[5996]<=26'd9733122; ROM4[5996]<=26'd23458213;
ROM1[5997]<=26'd1979419; ROM2[5997]<=26'd11139296; ROM3[5997]<=26'd9731430; ROM4[5997]<=26'd23459244;
ROM1[5998]<=26'd1997850; ROM2[5998]<=26'd11144451; ROM3[5998]<=26'd9734423; ROM4[5998]<=26'd23463086;
ROM1[5999]<=26'd2006939; ROM2[5999]<=26'd11146890; ROM3[5999]<=26'd9732508; ROM4[5999]<=26'd23463748;
ROM1[6000]<=26'd1996689; ROM2[6000]<=26'd11141385; ROM3[6000]<=26'd9729174; ROM4[6000]<=26'd23460227;
ROM1[6001]<=26'd1984752; ROM2[6001]<=26'd11136389; ROM3[6001]<=26'd9729929; ROM4[6001]<=26'd23457608;
ROM1[6002]<=26'd1981548; ROM2[6002]<=26'd11140445; ROM3[6002]<=26'd9738812; ROM4[6002]<=26'd23462694;
ROM1[6003]<=26'd1974881; ROM2[6003]<=26'd11138952; ROM3[6003]<=26'd9744094; ROM4[6003]<=26'd23462512;
ROM1[6004]<=26'd1968429; ROM2[6004]<=26'd11135123; ROM3[6004]<=26'd9741915; ROM4[6004]<=26'd23460162;
ROM1[6005]<=26'd1974771; ROM2[6005]<=26'd11137647; ROM3[6005]<=26'd9742877; ROM4[6005]<=26'd23461776;
ROM1[6006]<=26'd1989350; ROM2[6006]<=26'd11142096; ROM3[6006]<=26'd9741607; ROM4[6006]<=26'd23464301;
ROM1[6007]<=26'd2000566; ROM2[6007]<=26'd11145466; ROM3[6007]<=26'd9735527; ROM4[6007]<=26'd23465741;
ROM1[6008]<=26'd2000004; ROM2[6008]<=26'd11145467; ROM3[6008]<=26'd9734347; ROM4[6008]<=26'd23465529;
ROM1[6009]<=26'd1990794; ROM2[6009]<=26'd11143896; ROM3[6009]<=26'd9733648; ROM4[6009]<=26'd23464030;
ROM1[6010]<=26'd1984034; ROM2[6010]<=26'd11144308; ROM3[6010]<=26'd9736561; ROM4[6010]<=26'd23465800;
ROM1[6011]<=26'd1981049; ROM2[6011]<=26'd11145160; ROM3[6011]<=26'd9739783; ROM4[6011]<=26'd23467206;
ROM1[6012]<=26'd1976830; ROM2[6012]<=26'd11144578; ROM3[6012]<=26'd9742302; ROM4[6012]<=26'd23467525;
ROM1[6013]<=26'd1976321; ROM2[6013]<=26'd11143272; ROM3[6013]<=26'd9742624; ROM4[6013]<=26'd23466934;
ROM1[6014]<=26'd1985260; ROM2[6014]<=26'd11145433; ROM3[6014]<=26'd9740642; ROM4[6014]<=26'd23466476;
ROM1[6015]<=26'd1999291; ROM2[6015]<=26'd11148837; ROM3[6015]<=26'd9738333; ROM4[6015]<=26'd23468358;
ROM1[6016]<=26'd1997668; ROM2[6016]<=26'd11143174; ROM3[6016]<=26'd9733002; ROM4[6016]<=26'd23463815;
ROM1[6017]<=26'd1997019; ROM2[6017]<=26'd11146381; ROM3[6017]<=26'd9739978; ROM4[6017]<=26'd23466744;
ROM1[6018]<=26'd1993980; ROM2[6018]<=26'd11149204; ROM3[6018]<=26'd9746692; ROM4[6018]<=26'd23470032;
ROM1[6019]<=26'd1985429; ROM2[6019]<=26'd11145874; ROM3[6019]<=26'd9747103; ROM4[6019]<=26'd23466589;
ROM1[6020]<=26'd1978350; ROM2[6020]<=26'd11145434; ROM3[6020]<=26'd9748967; ROM4[6020]<=26'd23465565;
ROM1[6021]<=26'd1973922; ROM2[6021]<=26'd11141530; ROM3[6021]<=26'd9746511; ROM4[6021]<=26'd23461896;
ROM1[6022]<=26'd1974500; ROM2[6022]<=26'd11136725; ROM3[6022]<=26'd9740308; ROM4[6022]<=26'd23454750;
ROM1[6023]<=26'd1985096; ROM2[6023]<=26'd11134999; ROM3[6023]<=26'd9734785; ROM4[6023]<=26'd23454953;
ROM1[6024]<=26'd1996131; ROM2[6024]<=26'd11137938; ROM3[6024]<=26'd9736831; ROM4[6024]<=26'd23458717;
ROM1[6025]<=26'd1991147; ROM2[6025]<=26'd11137188; ROM3[6025]<=26'd9738091; ROM4[6025]<=26'd23457547;
ROM1[6026]<=26'd1985947; ROM2[6026]<=26'd11138961; ROM3[6026]<=26'd9743536; ROM4[6026]<=26'd23462611;
ROM1[6027]<=26'd1982608; ROM2[6027]<=26'd11139845; ROM3[6027]<=26'd9749595; ROM4[6027]<=26'd23463681;
ROM1[6028]<=26'd1970423; ROM2[6028]<=26'd11131305; ROM3[6028]<=26'd9744275; ROM4[6028]<=26'd23455558;
ROM1[6029]<=26'd1967646; ROM2[6029]<=26'd11130639; ROM3[6029]<=26'd9744923; ROM4[6029]<=26'd23456229;
ROM1[6030]<=26'd1974374; ROM2[6030]<=26'd11133104; ROM3[6030]<=26'd9745713; ROM4[6030]<=26'd23457963;
ROM1[6031]<=26'd1983154; ROM2[6031]<=26'd11133021; ROM3[6031]<=26'd9737722; ROM4[6031]<=26'd23455438;
ROM1[6032]<=26'd1995150; ROM2[6032]<=26'd11136938; ROM3[6032]<=26'd9734165; ROM4[6032]<=26'd23457671;
ROM1[6033]<=26'd1992705; ROM2[6033]<=26'd11137152; ROM3[6033]<=26'd9734035; ROM4[6033]<=26'd23457369;
ROM1[6034]<=26'd1980759; ROM2[6034]<=26'd11133873; ROM3[6034]<=26'd9733319; ROM4[6034]<=26'd23453508;
ROM1[6035]<=26'd1973975; ROM2[6035]<=26'd11133604; ROM3[6035]<=26'd9735334; ROM4[6035]<=26'd23452442;
ROM1[6036]<=26'd1971497; ROM2[6036]<=26'd11135528; ROM3[6036]<=26'd9739108; ROM4[6036]<=26'd23455912;
ROM1[6037]<=26'd1971682; ROM2[6037]<=26'd11140809; ROM3[6037]<=26'd9745474; ROM4[6037]<=26'd23461954;
ROM1[6038]<=26'd1974827; ROM2[6038]<=26'd11143490; ROM3[6038]<=26'd9747463; ROM4[6038]<=26'd23464758;
ROM1[6039]<=26'd1976065; ROM2[6039]<=26'd11136934; ROM3[6039]<=26'd9738901; ROM4[6039]<=26'd23459160;
ROM1[6040]<=26'd1987210; ROM2[6040]<=26'd11135445; ROM3[6040]<=26'd9732447; ROM4[6040]<=26'd23456246;
ROM1[6041]<=26'd1990288; ROM2[6041]<=26'd11136702; ROM3[6041]<=26'd9732180; ROM4[6041]<=26'd23457195;
ROM1[6042]<=26'd1987203; ROM2[6042]<=26'd11138858; ROM3[6042]<=26'd9736027; ROM4[6042]<=26'd23459688;
ROM1[6043]<=26'd1985317; ROM2[6043]<=26'd11144836; ROM3[6043]<=26'd9745027; ROM4[6043]<=26'd23467163;
ROM1[6044]<=26'd1979789; ROM2[6044]<=26'd11144967; ROM3[6044]<=26'd9750770; ROM4[6044]<=26'd23469389;
ROM1[6045]<=26'd1971113; ROM2[6045]<=26'd11139799; ROM3[6045]<=26'd9753575; ROM4[6045]<=26'd23467528;
ROM1[6046]<=26'd1965928; ROM2[6046]<=26'd11137198; ROM3[6046]<=26'd9753389; ROM4[6046]<=26'd23467488;
ROM1[6047]<=26'd1975221; ROM2[6047]<=26'd11140108; ROM3[6047]<=26'd9753994; ROM4[6047]<=26'd23469208;
ROM1[6048]<=26'd1991970; ROM2[6048]<=26'd11146780; ROM3[6048]<=26'd9753469; ROM4[6048]<=26'd23472085;
ROM1[6049]<=26'd2006812; ROM2[6049]<=26'd11156884; ROM3[6049]<=26'd9758309; ROM4[6049]<=26'd23479797;
ROM1[6050]<=26'd2004415; ROM2[6050]<=26'd11155997; ROM3[6050]<=26'd9761717; ROM4[6050]<=26'd23480847;
ROM1[6051]<=26'd1988872; ROM2[6051]<=26'd11146654; ROM3[6051]<=26'd9755177; ROM4[6051]<=26'd23472725;
ROM1[6052]<=26'd1981246; ROM2[6052]<=26'd11144653; ROM3[6052]<=26'd9756010; ROM4[6052]<=26'd23472739;
ROM1[6053]<=26'd1972917; ROM2[6053]<=26'd11141256; ROM3[6053]<=26'd9756443; ROM4[6053]<=26'd23470448;
ROM1[6054]<=26'd1965431; ROM2[6054]<=26'd11139322; ROM3[6054]<=26'd9753477; ROM4[6054]<=26'd23466813;
ROM1[6055]<=26'd1970545; ROM2[6055]<=26'd11143700; ROM3[6055]<=26'd9753276; ROM4[6055]<=26'd23468821;
ROM1[6056]<=26'd1985512; ROM2[6056]<=26'd11147395; ROM3[6056]<=26'd9752192; ROM4[6056]<=26'd23470680;
ROM1[6057]<=26'd1996461; ROM2[6057]<=26'd11147352; ROM3[6057]<=26'd9747145; ROM4[6057]<=26'd23471458;
ROM1[6058]<=26'd1998960; ROM2[6058]<=26'd11150922; ROM3[6058]<=26'd9748360; ROM4[6058]<=26'd23474159;
ROM1[6059]<=26'd1994577; ROM2[6059]<=26'd11153456; ROM3[6059]<=26'd9754274; ROM4[6059]<=26'd23476525;
ROM1[6060]<=26'd1984661; ROM2[6060]<=26'd11151226; ROM3[6060]<=26'd9753765; ROM4[6060]<=26'd23474216;
ROM1[6061]<=26'd1975363; ROM2[6061]<=26'd11148406; ROM3[6061]<=26'd9749420; ROM4[6061]<=26'd23471482;
ROM1[6062]<=26'd1969359; ROM2[6062]<=26'd11146610; ROM3[6062]<=26'd9748572; ROM4[6062]<=26'd23471088;
ROM1[6063]<=26'd1972125; ROM2[6063]<=26'd11147942; ROM3[6063]<=26'd9749680; ROM4[6063]<=26'd23472437;
ROM1[6064]<=26'd1981672; ROM2[6064]<=26'd11151355; ROM3[6064]<=26'd9747008; ROM4[6064]<=26'd23472167;
ROM1[6065]<=26'd1994238; ROM2[6065]<=26'd11151343; ROM3[6065]<=26'd9738452; ROM4[6065]<=26'd23468893;
ROM1[6066]<=26'd1995234; ROM2[6066]<=26'd11147516; ROM3[6066]<=26'd9734366; ROM4[6066]<=26'd23465610;
ROM1[6067]<=26'd1991127; ROM2[6067]<=26'd11148830; ROM3[6067]<=26'd9739502; ROM4[6067]<=26'd23467770;
ROM1[6068]<=26'd1983189; ROM2[6068]<=26'd11147626; ROM3[6068]<=26'd9743759; ROM4[6068]<=26'd23467491;
ROM1[6069]<=26'd1973586; ROM2[6069]<=26'd11142839; ROM3[6069]<=26'd9743752; ROM4[6069]<=26'd23463541;
ROM1[6070]<=26'd1971134; ROM2[6070]<=26'd11144674; ROM3[6070]<=26'd9748802; ROM4[6070]<=26'd23466085;
ROM1[6071]<=26'd1972479; ROM2[6071]<=26'd11147872; ROM3[6071]<=26'd9752400; ROM4[6071]<=26'd23468326;
ROM1[6072]<=26'd1980521; ROM2[6072]<=26'd11150221; ROM3[6072]<=26'd9753350; ROM4[6072]<=26'd23471730;
ROM1[6073]<=26'd1988622; ROM2[6073]<=26'd11147130; ROM3[6073]<=26'd9746813; ROM4[6073]<=26'd23468378;
ROM1[6074]<=26'd1989963; ROM2[6074]<=26'd11142013; ROM3[6074]<=26'd9741476; ROM4[6074]<=26'd23463523;
ROM1[6075]<=26'd1985865; ROM2[6075]<=26'd11140948; ROM3[6075]<=26'd9744428; ROM4[6075]<=26'd23463811;
ROM1[6076]<=26'd1982655; ROM2[6076]<=26'd11144696; ROM3[6076]<=26'd9751794; ROM4[6076]<=26'd23467115;
ROM1[6077]<=26'd1984673; ROM2[6077]<=26'd11152868; ROM3[6077]<=26'd9761717; ROM4[6077]<=26'd23474055;
ROM1[6078]<=26'd1972821; ROM2[6078]<=26'd11146673; ROM3[6078]<=26'd9757779; ROM4[6078]<=26'd23468342;
ROM1[6079]<=26'd1959946; ROM2[6079]<=26'd11136455; ROM3[6079]<=26'd9750988; ROM4[6079]<=26'd23460213;
ROM1[6080]<=26'd1961839; ROM2[6080]<=26'd11136406; ROM3[6080]<=26'd9748781; ROM4[6080]<=26'd23459534;
ROM1[6081]<=26'd1980006; ROM2[6081]<=26'd11145304; ROM3[6081]<=26'd9752528; ROM4[6081]<=26'd23465818;
ROM1[6082]<=26'd1997095; ROM2[6082]<=26'd11152703; ROM3[6082]<=26'd9752905; ROM4[6082]<=26'd23470807;
ROM1[6083]<=26'd1992366; ROM2[6083]<=26'd11147369; ROM3[6083]<=26'd9745670; ROM4[6083]<=26'd23466355;
ROM1[6084]<=26'd1983579; ROM2[6084]<=26'd11141653; ROM3[6084]<=26'd9743747; ROM4[6084]<=26'd23462896;
ROM1[6085]<=26'd1975687; ROM2[6085]<=26'd11137298; ROM3[6085]<=26'd9745380; ROM4[6085]<=26'd23460680;
ROM1[6086]<=26'd1971293; ROM2[6086]<=26'd11138626; ROM3[6086]<=26'd9747014; ROM4[6086]<=26'd23461430;
ROM1[6087]<=26'd1971634; ROM2[6087]<=26'd11145492; ROM3[6087]<=26'd9755438; ROM4[6087]<=26'd23467083;
ROM1[6088]<=26'd1968081; ROM2[6088]<=26'd11140944; ROM3[6088]<=26'd9751653; ROM4[6088]<=26'd23462326;
ROM1[6089]<=26'd1967835; ROM2[6089]<=26'd11133882; ROM3[6089]<=26'd9738044; ROM4[6089]<=26'd23454267;
ROM1[6090]<=26'd1986707; ROM2[6090]<=26'd11141518; ROM3[6090]<=26'd9741779; ROM4[6090]<=26'd23461386;
ROM1[6091]<=26'd1996527; ROM2[6091]<=26'd11148217; ROM3[6091]<=26'd9747998; ROM4[6091]<=26'd23467853;
ROM1[6092]<=26'd1990809; ROM2[6092]<=26'd11148459; ROM3[6092]<=26'd9749581; ROM4[6092]<=26'd23468571;
ROM1[6093]<=26'd1982096; ROM2[6093]<=26'd11145730; ROM3[6093]<=26'd9752007; ROM4[6093]<=26'd23468151;
ROM1[6094]<=26'd1974806; ROM2[6094]<=26'd11143499; ROM3[6094]<=26'd9752144; ROM4[6094]<=26'd23466512;
ROM1[6095]<=26'd1967316; ROM2[6095]<=26'd11140891; ROM3[6095]<=26'd9753240; ROM4[6095]<=26'd23465275;
ROM1[6096]<=26'd1965078; ROM2[6096]<=26'd11139851; ROM3[6096]<=26'd9753239; ROM4[6096]<=26'd23464243;
ROM1[6097]<=26'd1974726; ROM2[6097]<=26'd11145008; ROM3[6097]<=26'd9751971; ROM4[6097]<=26'd23466416;
ROM1[6098]<=26'd1985160; ROM2[6098]<=26'd11144180; ROM3[6098]<=26'd9743861; ROM4[6098]<=26'd23461928;
ROM1[6099]<=26'd1989024; ROM2[6099]<=26'd11140619; ROM3[6099]<=26'd9733235; ROM4[6099]<=26'd23456449;
ROM1[6100]<=26'd1984646; ROM2[6100]<=26'd11138956; ROM3[6100]<=26'd9732538; ROM4[6100]<=26'd23457096;
ROM1[6101]<=26'd1973545; ROM2[6101]<=26'd11134382; ROM3[6101]<=26'd9732733; ROM4[6101]<=26'd23454901;
ROM1[6102]<=26'd1968366; ROM2[6102]<=26'd11134917; ROM3[6102]<=26'd9735353; ROM4[6102]<=26'd23456738;
ROM1[6103]<=26'd1973557; ROM2[6103]<=26'd11145136; ROM3[6103]<=26'd9746776; ROM4[6103]<=26'd23466640;
ROM1[6104]<=26'd1971204; ROM2[6104]<=26'd11145422; ROM3[6104]<=26'd9748632; ROM4[6104]<=26'd23466533;
ROM1[6105]<=26'd1968944; ROM2[6105]<=26'd11139643; ROM3[6105]<=26'd9742406; ROM4[6105]<=26'd23460664;
ROM1[6106]<=26'd1975965; ROM2[6106]<=26'd11137290; ROM3[6106]<=26'd9737832; ROM4[6106]<=26'd23458331;
ROM1[6107]<=26'd1985833; ROM2[6107]<=26'd11137314; ROM3[6107]<=26'd9734415; ROM4[6107]<=26'd23457243;
ROM1[6108]<=26'd1988785; ROM2[6108]<=26'd11139160; ROM3[6108]<=26'd9736969; ROM4[6108]<=26'd23460666;
ROM1[6109]<=26'd1986897; ROM2[6109]<=26'd11143451; ROM3[6109]<=26'd9745948; ROM4[6109]<=26'd23467438;
ROM1[6110]<=26'd1984918; ROM2[6110]<=26'd11144444; ROM3[6110]<=26'd9753046; ROM4[6110]<=26'd23471174;
ROM1[6111]<=26'd1975119; ROM2[6111]<=26'd11138299; ROM3[6111]<=26'd9751612; ROM4[6111]<=26'd23468067;
ROM1[6112]<=26'd1965911; ROM2[6112]<=26'd11135504; ROM3[6112]<=26'd9751260; ROM4[6112]<=26'd23464913;
ROM1[6113]<=26'd1967173; ROM2[6113]<=26'd11135310; ROM3[6113]<=26'd9751706; ROM4[6113]<=26'd23462986;
ROM1[6114]<=26'd1974321; ROM2[6114]<=26'd11134652; ROM3[6114]<=26'd9746533; ROM4[6114]<=26'd23461901;
ROM1[6115]<=26'd1991167; ROM2[6115]<=26'd11140783; ROM3[6115]<=26'd9745045; ROM4[6115]<=26'd23467440;
ROM1[6116]<=26'd1995448; ROM2[6116]<=26'd11142959; ROM3[6116]<=26'd9744502; ROM4[6116]<=26'd23468786;
ROM1[6117]<=26'd1986939; ROM2[6117]<=26'd11141180; ROM3[6117]<=26'd9744501; ROM4[6117]<=26'd23467211;
ROM1[6118]<=26'd1982415; ROM2[6118]<=26'd11143461; ROM3[6118]<=26'd9750376; ROM4[6118]<=26'd23469315;
ROM1[6119]<=26'd1977777; ROM2[6119]<=26'd11142867; ROM3[6119]<=26'd9753277; ROM4[6119]<=26'd23468146;
ROM1[6120]<=26'd1976233; ROM2[6120]<=26'd11148572; ROM3[6120]<=26'd9760263; ROM4[6120]<=26'd23473792;
ROM1[6121]<=26'd1971238; ROM2[6121]<=26'd11146378; ROM3[6121]<=26'd9757328; ROM4[6121]<=26'd23470339;
ROM1[6122]<=26'd1967967; ROM2[6122]<=26'd11137753; ROM3[6122]<=26'd9744127; ROM4[6122]<=26'd23458766;
ROM1[6123]<=26'd1978945; ROM2[6123]<=26'd11137640; ROM3[6123]<=26'd9737443; ROM4[6123]<=26'd23458229;
ROM1[6124]<=26'd1985600; ROM2[6124]<=26'd11136699; ROM3[6124]<=26'd9734219; ROM4[6124]<=26'd23457477;
ROM1[6125]<=26'd1985036; ROM2[6125]<=26'd11138751; ROM3[6125]<=26'd9737080; ROM4[6125]<=26'd23458294;
ROM1[6126]<=26'd1980089; ROM2[6126]<=26'd11139996; ROM3[6126]<=26'd9741755; ROM4[6126]<=26'd23460327;
ROM1[6127]<=26'd1971803; ROM2[6127]<=26'd11136437; ROM3[6127]<=26'd9740958; ROM4[6127]<=26'd23457966;
ROM1[6128]<=26'd1963208; ROM2[6128]<=26'd11133739; ROM3[6128]<=26'd9737848; ROM4[6128]<=26'd23454960;
ROM1[6129]<=26'd1963405; ROM2[6129]<=26'd11135556; ROM3[6129]<=26'd9740078; ROM4[6129]<=26'd23457120;
ROM1[6130]<=26'd1970570; ROM2[6130]<=26'd11139620; ROM3[6130]<=26'd9741252; ROM4[6130]<=26'd23461134;
ROM1[6131]<=26'd1981253; ROM2[6131]<=26'd11142355; ROM3[6131]<=26'd9735866; ROM4[6131]<=26'd23459803;
ROM1[6132]<=26'd1992323; ROM2[6132]<=26'd11141534; ROM3[6132]<=26'd9730698; ROM4[6132]<=26'd23457328;
ROM1[6133]<=26'd1988475; ROM2[6133]<=26'd11138405; ROM3[6133]<=26'd9727779; ROM4[6133]<=26'd23456731;
ROM1[6134]<=26'd1989173; ROM2[6134]<=26'd11146350; ROM3[6134]<=26'd9736738; ROM4[6134]<=26'd23464250;
ROM1[6135]<=26'd1985913; ROM2[6135]<=26'd11148544; ROM3[6135]<=26'd9743103; ROM4[6135]<=26'd23468280;
ROM1[6136]<=26'd1973945; ROM2[6136]<=26'd11141209; ROM3[6136]<=26'd9736453; ROM4[6136]<=26'd23462178;
ROM1[6137]<=26'd1972047; ROM2[6137]<=26'd11143393; ROM3[6137]<=26'd9741079; ROM4[6137]<=26'd23465171;
ROM1[6138]<=26'd1971422; ROM2[6138]<=26'd11142754; ROM3[6138]<=26'd9741613; ROM4[6138]<=26'd23465512;
ROM1[6139]<=26'd1971512; ROM2[6139]<=26'd11137164; ROM3[6139]<=26'd9729779; ROM4[6139]<=26'd23456478;
ROM1[6140]<=26'd1983760; ROM2[6140]<=26'd11139163; ROM3[6140]<=26'd9725708; ROM4[6140]<=26'd23454205;
ROM1[6141]<=26'd1988121; ROM2[6141]<=26'd11140818; ROM3[6141]<=26'd9725585; ROM4[6141]<=26'd23454224;
ROM1[6142]<=26'd1981320; ROM2[6142]<=26'd11138118; ROM3[6142]<=26'd9725953; ROM4[6142]<=26'd23453400;
ROM1[6143]<=26'd1975433; ROM2[6143]<=26'd11137297; ROM3[6143]<=26'd9731070; ROM4[6143]<=26'd23454836;
ROM1[6144]<=26'd1971269; ROM2[6144]<=26'd11138542; ROM3[6144]<=26'd9734877; ROM4[6144]<=26'd23457198;
ROM1[6145]<=26'd1965693; ROM2[6145]<=26'd11139945; ROM3[6145]<=26'd9739040; ROM4[6145]<=26'd23459549;
ROM1[6146]<=26'd1967342; ROM2[6146]<=26'd11142561; ROM3[6146]<=26'd9741909; ROM4[6146]<=26'd23461638;
ROM1[6147]<=26'd1977760; ROM2[6147]<=26'd11145684; ROM3[6147]<=26'd9742759; ROM4[6147]<=26'd23463503;
ROM1[6148]<=26'd1987306; ROM2[6148]<=26'd11143160; ROM3[6148]<=26'd9737607; ROM4[6148]<=26'd23461262;
ROM1[6149]<=26'd1988203; ROM2[6149]<=26'd11136077; ROM3[6149]<=26'd9728715; ROM4[6149]<=26'd23455112;
ROM1[6150]<=26'd1979263; ROM2[6150]<=26'd11131485; ROM3[6150]<=26'd9728003; ROM4[6150]<=26'd23451175;
ROM1[6151]<=26'd1972021; ROM2[6151]<=26'd11130962; ROM3[6151]<=26'd9732833; ROM4[6151]<=26'd23452143;
ROM1[6152]<=26'd1972951; ROM2[6152]<=26'd11135252; ROM3[6152]<=26'd9742580; ROM4[6152]<=26'd23459113;
ROM1[6153]<=26'd1970592; ROM2[6153]<=26'd11138072; ROM3[6153]<=26'd9748259; ROM4[6153]<=26'd23462992;
ROM1[6154]<=26'd1967315; ROM2[6154]<=26'd11137139; ROM3[6154]<=26'd9748839; ROM4[6154]<=26'd23462462;
ROM1[6155]<=26'd1970542; ROM2[6155]<=26'd11137906; ROM3[6155]<=26'd9748834; ROM4[6155]<=26'd23463336;
ROM1[6156]<=26'd1981187; ROM2[6156]<=26'd11140456; ROM3[6156]<=26'd9743832; ROM4[6156]<=26'd23462882;
ROM1[6157]<=26'd1998266; ROM2[6157]<=26'd11148077; ROM3[6157]<=26'd9744822; ROM4[6157]<=26'd23469405;
ROM1[6158]<=26'd1997363; ROM2[6158]<=26'd11145825; ROM3[6158]<=26'd9742420; ROM4[6158]<=26'd23466770;
ROM1[6159]<=26'd1981921; ROM2[6159]<=26'd11134573; ROM3[6159]<=26'd9735086; ROM4[6159]<=26'd23457777;
ROM1[6160]<=26'd1977562; ROM2[6160]<=26'd11136158; ROM3[6160]<=26'd9740309; ROM4[6160]<=26'd23461392;
ROM1[6161]<=26'd1974543; ROM2[6161]<=26'd11138274; ROM3[6161]<=26'd9745089; ROM4[6161]<=26'd23463970;
ROM1[6162]<=26'd1969954; ROM2[6162]<=26'd11138850; ROM3[6162]<=26'd9747843; ROM4[6162]<=26'd23465883;
ROM1[6163]<=26'd1972667; ROM2[6163]<=26'd11140785; ROM3[6163]<=26'd9750390; ROM4[6163]<=26'd23467609;
ROM1[6164]<=26'd1977291; ROM2[6164]<=26'd11136562; ROM3[6164]<=26'd9744042; ROM4[6164]<=26'd23462381;
ROM1[6165]<=26'd1986055; ROM2[6165]<=26'd11133958; ROM3[6165]<=26'd9736057; ROM4[6165]<=26'd23459078;
ROM1[6166]<=26'd1989702; ROM2[6166]<=26'd11134564; ROM3[6166]<=26'd9736696; ROM4[6166]<=26'd23460454;
ROM1[6167]<=26'd1988733; ROM2[6167]<=26'd11139567; ROM3[6167]<=26'd9744569; ROM4[6167]<=26'd23465022;
ROM1[6168]<=26'd1987951; ROM2[6168]<=26'd11145203; ROM3[6168]<=26'd9754704; ROM4[6168]<=26'd23472002;
ROM1[6169]<=26'd1982254; ROM2[6169]<=26'd11142492; ROM3[6169]<=26'd9756125; ROM4[6169]<=26'd23469793;
ROM1[6170]<=26'd1968033; ROM2[6170]<=26'd11134530; ROM3[6170]<=26'd9749741; ROM4[6170]<=26'd23462101;
ROM1[6171]<=26'd1963616; ROM2[6171]<=26'd11131313; ROM3[6171]<=26'd9744777; ROM4[6171]<=26'd23458690;
ROM1[6172]<=26'd1968431; ROM2[6172]<=26'd11131544; ROM3[6172]<=26'd9741002; ROM4[6172]<=26'd23456424;
ROM1[6173]<=26'd1984789; ROM2[6173]<=26'd11136559; ROM3[6173]<=26'd9741897; ROM4[6173]<=26'd23461188;
ROM1[6174]<=26'd2002235; ROM2[6174]<=26'd11148021; ROM3[6174]<=26'd9750072; ROM4[6174]<=26'd23471530;
ROM1[6175]<=26'd1999102; ROM2[6175]<=26'd11150375; ROM3[6175]<=26'd9754095; ROM4[6175]<=26'd23474010;
ROM1[6176]<=26'd1987212; ROM2[6176]<=26'd11144588; ROM3[6176]<=26'd9753108; ROM4[6176]<=26'd23470808;
ROM1[6177]<=26'd1977701; ROM2[6177]<=26'd11140713; ROM3[6177]<=26'd9750550; ROM4[6177]<=26'd23465763;
ROM1[6178]<=26'd1966484; ROM2[6178]<=26'd11133704; ROM3[6178]<=26'd9746216; ROM4[6178]<=26'd23460251;
ROM1[6179]<=26'd1963616; ROM2[6179]<=26'd11131100; ROM3[6179]<=26'd9746153; ROM4[6179]<=26'd23458695;
ROM1[6180]<=26'd1970543; ROM2[6180]<=26'd11135211; ROM3[6180]<=26'd9746315; ROM4[6180]<=26'd23459851;
ROM1[6181]<=26'd1981517; ROM2[6181]<=26'd11137068; ROM3[6181]<=26'd9741441; ROM4[6181]<=26'd23460349;
ROM1[6182]<=26'd1988554; ROM2[6182]<=26'd11133284; ROM3[6182]<=26'd9732325; ROM4[6182]<=26'd23455024;
ROM1[6183]<=26'd1987464; ROM2[6183]<=26'd11133855; ROM3[6183]<=26'd9731841; ROM4[6183]<=26'd23454728;
ROM1[6184]<=26'd1982567; ROM2[6184]<=26'd11135825; ROM3[6184]<=26'd9737903; ROM4[6184]<=26'd23457982;
ROM1[6185]<=26'd1976672; ROM2[6185]<=26'd11135390; ROM3[6185]<=26'd9744190; ROM4[6185]<=26'd23459358;
ROM1[6186]<=26'd1972142; ROM2[6186]<=26'd11137575; ROM3[6186]<=26'd9747445; ROM4[6186]<=26'd23461693;
ROM1[6187]<=26'd1967319; ROM2[6187]<=26'd11136627; ROM3[6187]<=26'd9748285; ROM4[6187]<=26'd23462389;
ROM1[6188]<=26'd1970547; ROM2[6188]<=26'd11137177; ROM3[6188]<=26'd9747290; ROM4[6188]<=26'd23462415;
ROM1[6189]<=26'd1979202; ROM2[6189]<=26'd11138807; ROM3[6189]<=26'd9741061; ROM4[6189]<=26'd23460931;
ROM1[6190]<=26'd1991483; ROM2[6190]<=26'd11138727; ROM3[6190]<=26'd9734960; ROM4[6190]<=26'd23460182;
ROM1[6191]<=26'd1994409; ROM2[6191]<=26'd11139173; ROM3[6191]<=26'd9733216; ROM4[6191]<=26'd23460775;
ROM1[6192]<=26'd1986620; ROM2[6192]<=26'd11138277; ROM3[6192]<=26'd9733180; ROM4[6192]<=26'd23459353;
ROM1[6193]<=26'd1979660; ROM2[6193]<=26'd11138535; ROM3[6193]<=26'd9737427; ROM4[6193]<=26'd23459221;
ROM1[6194]<=26'd1971236; ROM2[6194]<=26'd11134836; ROM3[6194]<=26'd9737408; ROM4[6194]<=26'd23456506;
ROM1[6195]<=26'd1964955; ROM2[6195]<=26'd11133266; ROM3[6195]<=26'd9738889; ROM4[6195]<=26'd23454396;
ROM1[6196]<=26'd1964705; ROM2[6196]<=26'd11135361; ROM3[6196]<=26'd9741985; ROM4[6196]<=26'd23455846;
ROM1[6197]<=26'd1971461; ROM2[6197]<=26'd11135429; ROM3[6197]<=26'd9740427; ROM4[6197]<=26'd23456266;
ROM1[6198]<=26'd1988815; ROM2[6198]<=26'd11142550; ROM3[6198]<=26'd9740343; ROM4[6198]<=26'd23459869;
ROM1[6199]<=26'd1998569; ROM2[6199]<=26'd11147533; ROM3[6199]<=26'd9742397; ROM4[6199]<=26'd23463888;
ROM1[6200]<=26'd1993669; ROM2[6200]<=26'd11144399; ROM3[6200]<=26'd9743650; ROM4[6200]<=26'd23462763;
ROM1[6201]<=26'd1979836; ROM2[6201]<=26'd11136701; ROM3[6201]<=26'd9740610; ROM4[6201]<=26'd23456897;
ROM1[6202]<=26'd1971974; ROM2[6202]<=26'd11133010; ROM3[6202]<=26'd9743351; ROM4[6202]<=26'd23455976;
ROM1[6203]<=26'd1967625; ROM2[6203]<=26'd11133075; ROM3[6203]<=26'd9747735; ROM4[6203]<=26'd23457124;
ROM1[6204]<=26'd1966496; ROM2[6204]<=26'd11135754; ROM3[6204]<=26'd9750218; ROM4[6204]<=26'd23459986;
ROM1[6205]<=26'd1972635; ROM2[6205]<=26'd11139192; ROM3[6205]<=26'd9751149; ROM4[6205]<=26'd23461837;
ROM1[6206]<=26'd1987063; ROM2[6206]<=26'd11144080; ROM3[6206]<=26'd9747454; ROM4[6206]<=26'd23463109;
ROM1[6207]<=26'd1998047; ROM2[6207]<=26'd11145584; ROM3[6207]<=26'd9739565; ROM4[6207]<=26'd23462947;
ROM1[6208]<=26'd2001357; ROM2[6208]<=26'd11149114; ROM3[6208]<=26'd9742066; ROM4[6208]<=26'd23465803;
ROM1[6209]<=26'd1996247; ROM2[6209]<=26'd11150089; ROM3[6209]<=26'd9746312; ROM4[6209]<=26'd23468537;
ROM1[6210]<=26'd1979987; ROM2[6210]<=26'd11140647; ROM3[6210]<=26'd9742228; ROM4[6210]<=26'd23461868;
ROM1[6211]<=26'd1970237; ROM2[6211]<=26'd11134850; ROM3[6211]<=26'd9741098; ROM4[6211]<=26'd23457443;
ROM1[6212]<=26'd1966151; ROM2[6212]<=26'd11135674; ROM3[6212]<=26'd9743294; ROM4[6212]<=26'd23459192;
ROM1[6213]<=26'd1974288; ROM2[6213]<=26'd11143202; ROM3[6213]<=26'd9748024; ROM4[6213]<=26'd23464926;
ROM1[6214]<=26'd1989642; ROM2[6214]<=26'd11148511; ROM3[6214]<=26'd9750321; ROM4[6214]<=26'd23469203;
ROM1[6215]<=26'd2000356; ROM2[6215]<=26'd11147679; ROM3[6215]<=26'd9742939; ROM4[6215]<=26'd23467201;
ROM1[6216]<=26'd2001898; ROM2[6216]<=26'd11147055; ROM3[6216]<=26'd9742003; ROM4[6216]<=26'd23466984;
ROM1[6217]<=26'd1992780; ROM2[6217]<=26'd11144012; ROM3[6217]<=26'd9743668; ROM4[6217]<=26'd23465833;
ROM1[6218]<=26'd1981161; ROM2[6218]<=26'd11139541; ROM3[6218]<=26'd9744211; ROM4[6218]<=26'd23463090;
ROM1[6219]<=26'd1977930; ROM2[6219]<=26'd11140631; ROM3[6219]<=26'd9750196; ROM4[6219]<=26'd23466075;
ROM1[6220]<=26'd1974566; ROM2[6220]<=26'd11142171; ROM3[6220]<=26'd9752166; ROM4[6220]<=26'd23466245;
ROM1[6221]<=26'd1973544; ROM2[6221]<=26'd11141920; ROM3[6221]<=26'd9748780; ROM4[6221]<=26'd23463435;
ROM1[6222]<=26'd1975656; ROM2[6222]<=26'd11140092; ROM3[6222]<=26'd9740278; ROM4[6222]<=26'd23458878;
ROM1[6223]<=26'd1990241; ROM2[6223]<=26'd11144702; ROM3[6223]<=26'd9735855; ROM4[6223]<=26'd23460409;
ROM1[6224]<=26'd1991508; ROM2[6224]<=26'd11139336; ROM3[6224]<=26'd9728174; ROM4[6224]<=26'd23454564;
ROM1[6225]<=26'd1976552; ROM2[6225]<=26'd11126815; ROM3[6225]<=26'd9718642; ROM4[6225]<=26'd23443419;
ROM1[6226]<=26'd1973643; ROM2[6226]<=26'd11127736; ROM3[6226]<=26'd9724956; ROM4[6226]<=26'd23447357;
ROM1[6227]<=26'd1969388; ROM2[6227]<=26'd11129348; ROM3[6227]<=26'd9729294; ROM4[6227]<=26'd23449053;
ROM1[6228]<=26'd1962993; ROM2[6228]<=26'd11129896; ROM3[6228]<=26'd9730703; ROM4[6228]<=26'd23449959;
ROM1[6229]<=26'd1963947; ROM2[6229]<=26'd11132921; ROM3[6229]<=26'd9735680; ROM4[6229]<=26'd23452773;
ROM1[6230]<=26'd1968753; ROM2[6230]<=26'd11132702; ROM3[6230]<=26'd9735197; ROM4[6230]<=26'd23451507;
ROM1[6231]<=26'd1978070; ROM2[6231]<=26'd11130486; ROM3[6231]<=26'd9729198; ROM4[6231]<=26'd23449474;
ROM1[6232]<=26'd1984210; ROM2[6232]<=26'd11127157; ROM3[6232]<=26'd9721305; ROM4[6232]<=26'd23446414;
ROM1[6233]<=26'd1984824; ROM2[6233]<=26'd11129026; ROM3[6233]<=26'd9723802; ROM4[6233]<=26'd23450646;
ROM1[6234]<=26'd1987312; ROM2[6234]<=26'd11136478; ROM3[6234]<=26'd9733448; ROM4[6234]<=26'd23459073;
ROM1[6235]<=26'd1981040; ROM2[6235]<=26'd11136523; ROM3[6235]<=26'd9737196; ROM4[6235]<=26'd23459422;
ROM1[6236]<=26'd1973949; ROM2[6236]<=26'd11132708; ROM3[6236]<=26'd9736443; ROM4[6236]<=26'd23458178;
ROM1[6237]<=26'd1974466; ROM2[6237]<=26'd11137149; ROM3[6237]<=26'd9743944; ROM4[6237]<=26'd23463109;
ROM1[6238]<=26'd1975113; ROM2[6238]<=26'd11139351; ROM3[6238]<=26'd9744151; ROM4[6238]<=26'd23462645;
ROM1[6239]<=26'd1973799; ROM2[6239]<=26'd11131211; ROM3[6239]<=26'd9730681; ROM4[6239]<=26'd23452469;
ROM1[6240]<=26'd1981444; ROM2[6240]<=26'd11126934; ROM3[6240]<=26'd9721744; ROM4[6240]<=26'd23447088;
ROM1[6241]<=26'd1982375; ROM2[6241]<=26'd11124533; ROM3[6241]<=26'd9719625; ROM4[6241]<=26'd23445240;
ROM1[6242]<=26'd1972590; ROM2[6242]<=26'd11120875; ROM3[6242]<=26'd9720414; ROM4[6242]<=26'd23442437;
ROM1[6243]<=26'd1968401; ROM2[6243]<=26'd11123448; ROM3[6243]<=26'd9728277; ROM4[6243]<=26'd23447672;
ROM1[6244]<=26'd1966747; ROM2[6244]<=26'd11126801; ROM3[6244]<=26'd9734965; ROM4[6244]<=26'd23452583;
ROM1[6245]<=26'd1959729; ROM2[6245]<=26'd11126295; ROM3[6245]<=26'd9736185; ROM4[6245]<=26'd23450690;
ROM1[6246]<=26'd1962873; ROM2[6246]<=26'd11129812; ROM3[6246]<=26'd9740750; ROM4[6246]<=26'd23454600;
ROM1[6247]<=26'd1974120; ROM2[6247]<=26'd11133731; ROM3[6247]<=26'd9741432; ROM4[6247]<=26'd23456385;
ROM1[6248]<=26'd1989369; ROM2[6248]<=26'd11137542; ROM3[6248]<=26'd9738642; ROM4[6248]<=26'd23456472;
ROM1[6249]<=26'd1996703; ROM2[6249]<=26'd11139446; ROM3[6249]<=26'd9737478; ROM4[6249]<=26'd23459283;
ROM1[6250]<=26'd1985316; ROM2[6250]<=26'd11131334; ROM3[6250]<=26'd9731431; ROM4[6250]<=26'd23453245;
ROM1[6251]<=26'd1977953; ROM2[6251]<=26'd11129726; ROM3[6251]<=26'd9734390; ROM4[6251]<=26'd23452652;
ROM1[6252]<=26'd1972652; ROM2[6252]<=26'd11130257; ROM3[6252]<=26'd9738222; ROM4[6252]<=26'd23454725;
ROM1[6253]<=26'd1966733; ROM2[6253]<=26'd11130930; ROM3[6253]<=26'd9738605; ROM4[6253]<=26'd23455104;
ROM1[6254]<=26'd1970004; ROM2[6254]<=26'd11139683; ROM3[6254]<=26'd9744191; ROM4[6254]<=26'd23460757;
ROM1[6255]<=26'd1977068; ROM2[6255]<=26'd11142592; ROM3[6255]<=26'd9744717; ROM4[6255]<=26'd23462427;
ROM1[6256]<=26'd1987192; ROM2[6256]<=26'd11141520; ROM3[6256]<=26'd9739887; ROM4[6256]<=26'd23460406;
ROM1[6257]<=26'd1995606; ROM2[6257]<=26'd11140878; ROM3[6257]<=26'd9733430; ROM4[6257]<=26'd23460731;
ROM1[6258]<=26'd1994671; ROM2[6258]<=26'd11140792; ROM3[6258]<=26'd9734708; ROM4[6258]<=26'd23462578;
ROM1[6259]<=26'd1986418; ROM2[6259]<=26'd11139530; ROM3[6259]<=26'd9737834; ROM4[6259]<=26'd23463419;
ROM1[6260]<=26'd1978751; ROM2[6260]<=26'd11138404; ROM3[6260]<=26'd9739104; ROM4[6260]<=26'd23462371;
ROM1[6261]<=26'd1970042; ROM2[6261]<=26'd11135572; ROM3[6261]<=26'd9736503; ROM4[6261]<=26'd23456766;
ROM1[6262]<=26'd1965949; ROM2[6262]<=26'd11136818; ROM3[6262]<=26'd9738518; ROM4[6262]<=26'd23457854;
ROM1[6263]<=26'd1973737; ROM2[6263]<=26'd11145608; ROM3[6263]<=26'd9744794; ROM4[6263]<=26'd23464221;
ROM1[6264]<=26'd1977358; ROM2[6264]<=26'd11143307; ROM3[6264]<=26'd9736725; ROM4[6264]<=26'd23458895;
ROM1[6265]<=26'd1982963; ROM2[6265]<=26'd11137569; ROM3[6265]<=26'd9727472; ROM4[6265]<=26'd23452751;
ROM1[6266]<=26'd1983092; ROM2[6266]<=26'd11133619; ROM3[6266]<=26'd9725411; ROM4[6266]<=26'd23451734;
ROM1[6267]<=26'd1974914; ROM2[6267]<=26'd11130348; ROM3[6267]<=26'd9726331; ROM4[6267]<=26'd23451357;
ROM1[6268]<=26'd1972507; ROM2[6268]<=26'd11133944; ROM3[6268]<=26'd9733766; ROM4[6268]<=26'd23456645;
ROM1[6269]<=26'd1973424; ROM2[6269]<=26'd11137948; ROM3[6269]<=26'd9741037; ROM4[6269]<=26'd23461247;
ROM1[6270]<=26'd1965154; ROM2[6270]<=26'd11136615; ROM3[6270]<=26'd9740823; ROM4[6270]<=26'd23458927;
ROM1[6271]<=26'd1958532; ROM2[6271]<=26'd11131774; ROM3[6271]<=26'd9734067; ROM4[6271]<=26'd23453105;
ROM1[6272]<=26'd1967466; ROM2[6272]<=26'd11132159; ROM3[6272]<=26'd9733445; ROM4[6272]<=26'd23454518;
ROM1[6273]<=26'd1983938; ROM2[6273]<=26'd11136320; ROM3[6273]<=26'd9733325; ROM4[6273]<=26'd23458279;
ROM1[6274]<=26'd1991390; ROM2[6274]<=26'd11136472; ROM3[6274]<=26'd9730473; ROM4[6274]<=26'd23456149;
ROM1[6275]<=26'd1985360; ROM2[6275]<=26'd11133306; ROM3[6275]<=26'd9732087; ROM4[6275]<=26'd23454645;
ROM1[6276]<=26'd1983041; ROM2[6276]<=26'd11138221; ROM3[6276]<=26'd9740249; ROM4[6276]<=26'd23459000;
ROM1[6277]<=26'd1982868; ROM2[6277]<=26'd11142737; ROM3[6277]<=26'd9747372; ROM4[6277]<=26'd23464533;
ROM1[6278]<=26'd1967648; ROM2[6278]<=26'd11131276; ROM3[6278]<=26'd9739805; ROM4[6278]<=26'd23456582;
ROM1[6279]<=26'd1965037; ROM2[6279]<=26'd11131599; ROM3[6279]<=26'd9739915; ROM4[6279]<=26'd23456093;
ROM1[6280]<=26'd1972903; ROM2[6280]<=26'd11138416; ROM3[6280]<=26'd9742154; ROM4[6280]<=26'd23461398;
ROM1[6281]<=26'd1975518; ROM2[6281]<=26'd11133158; ROM3[6281]<=26'd9729303; ROM4[6281]<=26'd23453043;
ROM1[6282]<=26'd1984591; ROM2[6282]<=26'd11134062; ROM3[6282]<=26'd9722562; ROM4[6282]<=26'd23451893;
ROM1[6283]<=26'd1987294; ROM2[6283]<=26'd11137436; ROM3[6283]<=26'd9725365; ROM4[6283]<=26'd23456645;
ROM1[6284]<=26'd1981765; ROM2[6284]<=26'd11135217; ROM3[6284]<=26'd9728045; ROM4[6284]<=26'd23456781;
ROM1[6285]<=26'd1975838; ROM2[6285]<=26'd11134249; ROM3[6285]<=26'd9732175; ROM4[6285]<=26'd23457396;
ROM1[6286]<=26'd1975046; ROM2[6286]<=26'd11138951; ROM3[6286]<=26'd9739926; ROM4[6286]<=26'd23462904;
ROM1[6287]<=26'd1970482; ROM2[6287]<=26'd11139509; ROM3[6287]<=26'd9742326; ROM4[6287]<=26'd23464424;
ROM1[6288]<=26'd1970066; ROM2[6288]<=26'd11139389; ROM3[6288]<=26'd9742137; ROM4[6288]<=26'd23464269;
ROM1[6289]<=26'd1985353; ROM2[6289]<=26'd11146392; ROM3[6289]<=26'd9744399; ROM4[6289]<=26'd23469395;
ROM1[6290]<=26'd2002295; ROM2[6290]<=26'd11151780; ROM3[6290]<=26'd9745708; ROM4[6290]<=26'd23472875;
ROM1[6291]<=26'd2001968; ROM2[6291]<=26'd11151665; ROM3[6291]<=26'd9744746; ROM4[6291]<=26'd23471248;
ROM1[6292]<=26'd1990968; ROM2[6292]<=26'd11145907; ROM3[6292]<=26'd9740358; ROM4[6292]<=26'd23464092;
ROM1[6293]<=26'd1980499; ROM2[6293]<=26'd11139653; ROM3[6293]<=26'd9740015; ROM4[6293]<=26'd23460096;
ROM1[6294]<=26'd1974696; ROM2[6294]<=26'd11139516; ROM3[6294]<=26'd9744139; ROM4[6294]<=26'd23461544;
ROM1[6295]<=26'd1967991; ROM2[6295]<=26'd11137540; ROM3[6295]<=26'd9747733; ROM4[6295]<=26'd23461166;
ROM1[6296]<=26'd1968077; ROM2[6296]<=26'd11137905; ROM3[6296]<=26'd9750802; ROM4[6296]<=26'd23464713;
ROM1[6297]<=26'd1980912; ROM2[6297]<=26'd11146211; ROM3[6297]<=26'd9755338; ROM4[6297]<=26'd23471981;
ROM1[6298]<=26'd2004743; ROM2[6298]<=26'd11158624; ROM3[6298]<=26'd9757813; ROM4[6298]<=26'd23479905;
ROM1[6299]<=26'd2009314; ROM2[6299]<=26'd11156277; ROM3[6299]<=26'd9750093; ROM4[6299]<=26'd23476986;
ROM1[6300]<=26'd1996010; ROM2[6300]<=26'd11146836; ROM3[6300]<=26'd9744889; ROM4[6300]<=26'd23468366;
ROM1[6301]<=26'd1989898; ROM2[6301]<=26'd11150700; ROM3[6301]<=26'd9750605; ROM4[6301]<=26'd23470483;
ROM1[6302]<=26'd1983693; ROM2[6302]<=26'd11150221; ROM3[6302]<=26'd9752732; ROM4[6302]<=26'd23469832;
ROM1[6303]<=26'd1972490; ROM2[6303]<=26'd11142471; ROM3[6303]<=26'd9750969; ROM4[6303]<=26'd23464835;
ROM1[6304]<=26'd1967971; ROM2[6304]<=26'd11142735; ROM3[6304]<=26'd9752121; ROM4[6304]<=26'd23464301;
ROM1[6305]<=26'd1967406; ROM2[6305]<=26'd11138463; ROM3[6305]<=26'd9745573; ROM4[6305]<=26'd23458211;
ROM1[6306]<=26'd1973843; ROM2[6306]<=26'd11135242; ROM3[6306]<=26'd9737482; ROM4[6306]<=26'd23455040;
ROM1[6307]<=26'd1990425; ROM2[6307]<=26'd11144039; ROM3[6307]<=26'd9739352; ROM4[6307]<=26'd23461873;
ROM1[6308]<=26'd1993031; ROM2[6308]<=26'd11148123; ROM3[6308]<=26'd9743546; ROM4[6308]<=26'd23466535;
ROM1[6309]<=26'd1982469; ROM2[6309]<=26'd11144409; ROM3[6309]<=26'd9744447; ROM4[6309]<=26'd23466041;
ROM1[6310]<=26'd1978689; ROM2[6310]<=26'd11144954; ROM3[6310]<=26'd9750369; ROM4[6310]<=26'd23469944;
ROM1[6311]<=26'd1980173; ROM2[6311]<=26'd11152595; ROM3[6311]<=26'd9759034; ROM4[6311]<=26'd23475729;
ROM1[6312]<=26'd1970869; ROM2[6312]<=26'd11147418; ROM3[6312]<=26'd9754623; ROM4[6312]<=26'd23471062;
ROM1[6313]<=26'd1963719; ROM2[6313]<=26'd11136977; ROM3[6313]<=26'd9743404; ROM4[6313]<=26'd23461532;
ROM1[6314]<=26'd1965930; ROM2[6314]<=26'd11132146; ROM3[6314]<=26'd9733204; ROM4[6314]<=26'd23451707;
ROM1[6315]<=26'd1975730; ROM2[6315]<=26'd11129475; ROM3[6315]<=26'd9725123; ROM4[6315]<=26'd23448525;
ROM1[6316]<=26'd1980602; ROM2[6316]<=26'd11130433; ROM3[6316]<=26'd9725444; ROM4[6316]<=26'd23450690;
ROM1[6317]<=26'd1973875; ROM2[6317]<=26'd11130658; ROM3[6317]<=26'd9728994; ROM4[6317]<=26'd23453088;
ROM1[6318]<=26'd1963301; ROM2[6318]<=26'd11128318; ROM3[6318]<=26'd9732689; ROM4[6318]<=26'd23453685;
ROM1[6319]<=26'd1961683; ROM2[6319]<=26'd11129605; ROM3[6319]<=26'd9739805; ROM4[6319]<=26'd23456051;
ROM1[6320]<=26'd1961371; ROM2[6320]<=26'd11134361; ROM3[6320]<=26'd9746953; ROM4[6320]<=26'd23461176;
ROM1[6321]<=26'd1958278; ROM2[6321]<=26'd11133360; ROM3[6321]<=26'd9744984; ROM4[6321]<=26'd23459293;
ROM1[6322]<=26'd1962360; ROM2[6322]<=26'd11130976; ROM3[6322]<=26'd9739502; ROM4[6322]<=26'd23454957;
ROM1[6323]<=26'd1971947; ROM2[6323]<=26'd11129339; ROM3[6323]<=26'd9732313; ROM4[6323]<=26'd23452739;
ROM1[6324]<=26'd1976589; ROM2[6324]<=26'd11128869; ROM3[6324]<=26'd9729339; ROM4[6324]<=26'd23452141;
ROM1[6325]<=26'd1975561; ROM2[6325]<=26'd11131741; ROM3[6325]<=26'd9736244; ROM4[6325]<=26'd23454989;
ROM1[6326]<=26'd1972001; ROM2[6326]<=26'd11134133; ROM3[6326]<=26'd9743843; ROM4[6326]<=26'd23459942;
ROM1[6327]<=26'd1964938; ROM2[6327]<=26'd11131328; ROM3[6327]<=26'd9744996; ROM4[6327]<=26'd23457885;
ROM1[6328]<=26'd1961917; ROM2[6328]<=26'd11132343; ROM3[6328]<=26'd9747152; ROM4[6328]<=26'd23457997;
ROM1[6329]<=26'd1967512; ROM2[6329]<=26'd11138005; ROM3[6329]<=26'd9754256; ROM4[6329]<=26'd23464814;
ROM1[6330]<=26'd1967023; ROM2[6330]<=26'd11133748; ROM3[6330]<=26'd9747557; ROM4[6330]<=26'd23461067;
ROM1[6331]<=26'd1973080; ROM2[6331]<=26'd11131912; ROM3[6331]<=26'd9739943; ROM4[6331]<=26'd23458939;
ROM1[6332]<=26'd1981605; ROM2[6332]<=26'd11132287; ROM3[6332]<=26'd9735592; ROM4[6332]<=26'd23457762;
ROM1[6333]<=26'd1979539; ROM2[6333]<=26'd11131594; ROM3[6333]<=26'd9735279; ROM4[6333]<=26'd23457104;
ROM1[6334]<=26'd1977579; ROM2[6334]<=26'd11136503; ROM3[6334]<=26'd9742596; ROM4[6334]<=26'd23461873;
ROM1[6335]<=26'd1978834; ROM2[6335]<=26'd11143625; ROM3[6335]<=26'd9750878; ROM4[6335]<=26'd23468378;
ROM1[6336]<=26'd1980321; ROM2[6336]<=26'd11149930; ROM3[6336]<=26'd9759955; ROM4[6336]<=26'd23475579;
ROM1[6337]<=26'd1970962; ROM2[6337]<=26'd11143527; ROM3[6337]<=26'd9756706; ROM4[6337]<=26'd23469573;
ROM1[6338]<=26'd1967484; ROM2[6338]<=26'd11138193; ROM3[6338]<=26'd9749708; ROM4[6338]<=26'd23463632;
ROM1[6339]<=26'd1978596; ROM2[6339]<=26'd11140128; ROM3[6339]<=26'd9746614; ROM4[6339]<=26'd23465277;
ROM1[6340]<=26'd1990690; ROM2[6340]<=26'd11138307; ROM3[6340]<=26'd9739238; ROM4[6340]<=26'd23463446;
ROM1[6341]<=26'd1990397; ROM2[6341]<=26'd11137629; ROM3[6341]<=26'd9735487; ROM4[6341]<=26'd23461904;
ROM1[6342]<=26'd1984966; ROM2[6342]<=26'd11137170; ROM3[6342]<=26'd9738445; ROM4[6342]<=26'd23463421;
ROM1[6343]<=26'd1976710; ROM2[6343]<=26'd11135586; ROM3[6343]<=26'd9742393; ROM4[6343]<=26'd23461704;
ROM1[6344]<=26'd1967880; ROM2[6344]<=26'd11131830; ROM3[6344]<=26'd9743071; ROM4[6344]<=26'd23457450;
ROM1[6345]<=26'd1965743; ROM2[6345]<=26'd11131843; ROM3[6345]<=26'd9748397; ROM4[6345]<=26'd23459682;
ROM1[6346]<=26'd1973132; ROM2[6346]<=26'd11139557; ROM3[6346]<=26'd9756349; ROM4[6346]<=26'd23466911;
ROM1[6347]<=26'd1983643; ROM2[6347]<=26'd11144023; ROM3[6347]<=26'd9755534; ROM4[6347]<=26'd23470323;
ROM1[6348]<=26'd1987228; ROM2[6348]<=26'd11137266; ROM3[6348]<=26'd9741579; ROM4[6348]<=26'd23461836;
ROM1[6349]<=26'd1990554; ROM2[6349]<=26'd11136283; ROM3[6349]<=26'd9734345; ROM4[6349]<=26'd23457960;
ROM1[6350]<=26'd1989603; ROM2[6350]<=26'd11139285; ROM3[6350]<=26'd9739057; ROM4[6350]<=26'd23460367;
ROM1[6351]<=26'd1978814; ROM2[6351]<=26'd11134812; ROM3[6351]<=26'd9739629; ROM4[6351]<=26'd23456345;
ROM1[6352]<=26'd1973046; ROM2[6352]<=26'd11135365; ROM3[6352]<=26'd9743453; ROM4[6352]<=26'd23458257;
ROM1[6353]<=26'd1969406; ROM2[6353]<=26'd11137346; ROM3[6353]<=26'd9748962; ROM4[6353]<=26'd23462457;
ROM1[6354]<=26'd1966435; ROM2[6354]<=26'd11136321; ROM3[6354]<=26'd9748495; ROM4[6354]<=26'd23462501;
ROM1[6355]<=26'd1968761; ROM2[6355]<=26'd11135760; ROM3[6355]<=26'd9747297; ROM4[6355]<=26'd23462274;
ROM1[6356]<=26'd1978942; ROM2[6356]<=26'd11135540; ROM3[6356]<=26'd9740716; ROM4[6356]<=26'd23460616;
ROM1[6357]<=26'd1987506; ROM2[6357]<=26'd11134724; ROM3[6357]<=26'd9733746; ROM4[6357]<=26'd23459538;
ROM1[6358]<=26'd1980462; ROM2[6358]<=26'd11129848; ROM3[6358]<=26'd9730642; ROM4[6358]<=26'd23455685;
ROM1[6359]<=26'd1976631; ROM2[6359]<=26'd11131666; ROM3[6359]<=26'd9734835; ROM4[6359]<=26'd23458120;
ROM1[6360]<=26'd1981149; ROM2[6360]<=26'd11141856; ROM3[6360]<=26'd9749373; ROM4[6360]<=26'd23469549;
ROM1[6361]<=26'd1976995; ROM2[6361]<=26'd11140502; ROM3[6361]<=26'd9751857; ROM4[6361]<=26'd23469246;
ROM1[6362]<=26'd1971736; ROM2[6362]<=26'd11140058; ROM3[6362]<=26'd9752595; ROM4[6362]<=26'd23468373;
ROM1[6363]<=26'd1968376; ROM2[6363]<=26'd11136993; ROM3[6363]<=26'd9748735; ROM4[6363]<=26'd23465195;
ROM1[6364]<=26'd1971833; ROM2[6364]<=26'd11131743; ROM3[6364]<=26'd9741079; ROM4[6364]<=26'd23459870;
ROM1[6365]<=26'd1986715; ROM2[6365]<=26'd11135897; ROM3[6365]<=26'd9740539; ROM4[6365]<=26'd23462558;
ROM1[6366]<=26'd1988730; ROM2[6366]<=26'd11135710; ROM3[6366]<=26'd9739874; ROM4[6366]<=26'd23463352;
ROM1[6367]<=26'd1984063; ROM2[6367]<=26'd11136447; ROM3[6367]<=26'd9743866; ROM4[6367]<=26'd23465887;
ROM1[6368]<=26'd1980088; ROM2[6368]<=26'd11137490; ROM3[6368]<=26'd9750132; ROM4[6368]<=26'd23468437;
ROM1[6369]<=26'd1975154; ROM2[6369]<=26'd11137756; ROM3[6369]<=26'd9752711; ROM4[6369]<=26'd23468784;
ROM1[6370]<=26'd1969133; ROM2[6370]<=26'd11136999; ROM3[6370]<=26'd9752184; ROM4[6370]<=26'd23469267;
ROM1[6371]<=26'd1968129; ROM2[6371]<=26'd11136387; ROM3[6371]<=26'd9749834; ROM4[6371]<=26'd23467664;
ROM1[6372]<=26'd1974133; ROM2[6372]<=26'd11137615; ROM3[6372]<=26'd9743889; ROM4[6372]<=26'd23465042;
ROM1[6373]<=26'd1985715; ROM2[6373]<=26'd11140723; ROM3[6373]<=26'd9736927; ROM4[6373]<=26'd23465763;
ROM1[6374]<=26'd1996235; ROM2[6374]<=26'd11145339; ROM3[6374]<=26'd9739171; ROM4[6374]<=26'd23469167;
ROM1[6375]<=26'd1998330; ROM2[6375]<=26'd11151831; ROM3[6375]<=26'd9748294; ROM4[6375]<=26'd23475690;
ROM1[6376]<=26'd1999012; ROM2[6376]<=26'd11158893; ROM3[6376]<=26'd9759669; ROM4[6376]<=26'd23485029;
ROM1[6377]<=26'd1993161; ROM2[6377]<=26'd11155699; ROM3[6377]<=26'd9762781; ROM4[6377]<=26'd23484055;
ROM1[6378]<=26'd1974950; ROM2[6378]<=26'd11143748; ROM3[6378]<=26'd9755317; ROM4[6378]<=26'd23473149;
ROM1[6379]<=26'd1964894; ROM2[6379]<=26'd11134693; ROM3[6379]<=26'd9750183; ROM4[6379]<=26'd23466712;
ROM1[6380]<=26'd1966653; ROM2[6380]<=26'd11133012; ROM3[6380]<=26'd9748327; ROM4[6380]<=26'd23465779;
ROM1[6381]<=26'd1979400; ROM2[6381]<=26'd11136523; ROM3[6381]<=26'd9747314; ROM4[6381]<=26'd23467899;
ROM1[6382]<=26'd1995994; ROM2[6382]<=26'd11142496; ROM3[6382]<=26'd9749164; ROM4[6382]<=26'd23471312;
ROM1[6383]<=26'd1993199; ROM2[6383]<=26'd11140702; ROM3[6383]<=26'd9746887; ROM4[6383]<=26'd23468614;
ROM1[6384]<=26'd1981891; ROM2[6384]<=26'd11135237; ROM3[6384]<=26'd9745612; ROM4[6384]<=26'd23464739;
ROM1[6385]<=26'd1977908; ROM2[6385]<=26'd11137706; ROM3[6385]<=26'd9752950; ROM4[6385]<=26'd23467962;
ROM1[6386]<=26'd1977434; ROM2[6386]<=26'd11141246; ROM3[6386]<=26'd9759692; ROM4[6386]<=26'd23474301;
ROM1[6387]<=26'd1969761; ROM2[6387]<=26'd11137475; ROM3[6387]<=26'd9759457; ROM4[6387]<=26'd23472083;
ROM1[6388]<=26'd1971942; ROM2[6388]<=26'd11139322; ROM3[6388]<=26'd9760650; ROM4[6388]<=26'd23472051;
ROM1[6389]<=26'd1980631; ROM2[6389]<=26'd11140694; ROM3[6389]<=26'd9757268; ROM4[6389]<=26'd23471846;
ROM1[6390]<=26'd1985525; ROM2[6390]<=26'd11135735; ROM3[6390]<=26'd9745723; ROM4[6390]<=26'd23464953;
ROM1[6391]<=26'd1987986; ROM2[6391]<=26'd11137416; ROM3[6391]<=26'd9744776; ROM4[6391]<=26'd23465262;
ROM1[6392]<=26'd1978992; ROM2[6392]<=26'd11135318; ROM3[6392]<=26'd9743779; ROM4[6392]<=26'd23462017;
ROM1[6393]<=26'd1967329; ROM2[6393]<=26'd11130400; ROM3[6393]<=26'd9742362; ROM4[6393]<=26'd23457790;
ROM1[6394]<=26'd1962766; ROM2[6394]<=26'd11130572; ROM3[6394]<=26'd9744751; ROM4[6394]<=26'd23459811;
ROM1[6395]<=26'd1954867; ROM2[6395]<=26'd11129038; ROM3[6395]<=26'd9745614; ROM4[6395]<=26'd23456723;
ROM1[6396]<=26'd1950876; ROM2[6396]<=26'd11127034; ROM3[6396]<=26'd9744904; ROM4[6396]<=26'd23454952;
ROM1[6397]<=26'd1958945; ROM2[6397]<=26'd11128795; ROM3[6397]<=26'd9741952; ROM4[6397]<=26'd23454670;
ROM1[6398]<=26'd1975267; ROM2[6398]<=26'd11133769; ROM3[6398]<=26'd9738988; ROM4[6398]<=26'd23456048;
ROM1[6399]<=26'd1984965; ROM2[6399]<=26'd11138363; ROM3[6399]<=26'd9738704; ROM4[6399]<=26'd23461917;
ROM1[6400]<=26'd1986910; ROM2[6400]<=26'd11144666; ROM3[6400]<=26'd9745288; ROM4[6400]<=26'd23467733;
ROM1[6401]<=26'd1980068; ROM2[6401]<=26'd11145762; ROM3[6401]<=26'd9750750; ROM4[6401]<=26'd23470624;
ROM1[6402]<=26'd1967228; ROM2[6402]<=26'd11138763; ROM3[6402]<=26'd9748295; ROM4[6402]<=26'd23465010;
ROM1[6403]<=26'd1960754; ROM2[6403]<=26'd11136892; ROM3[6403]<=26'd9752034; ROM4[6403]<=26'd23463469;
ROM1[6404]<=26'd1957021; ROM2[6404]<=26'd11134927; ROM3[6404]<=26'd9752314; ROM4[6404]<=26'd23463567;
ROM1[6405]<=26'd1959446; ROM2[6405]<=26'd11131502; ROM3[6405]<=26'd9746133; ROM4[6405]<=26'd23459862;
ROM1[6406]<=26'd1965094; ROM2[6406]<=26'd11129521; ROM3[6406]<=26'd9736565; ROM4[6406]<=26'd23454253;
ROM1[6407]<=26'd1972643; ROM2[6407]<=26'd11129948; ROM3[6407]<=26'd9728364; ROM4[6407]<=26'd23452202;
ROM1[6408]<=26'd1968897; ROM2[6408]<=26'd11127647; ROM3[6408]<=26'd9726198; ROM4[6408]<=26'd23450504;
ROM1[6409]<=26'd1962603; ROM2[6409]<=26'd11127790; ROM3[6409]<=26'd9729731; ROM4[6409]<=26'd23451329;
ROM1[6410]<=26'd1959633; ROM2[6410]<=26'd11128692; ROM3[6410]<=26'd9734342; ROM4[6410]<=26'd23451999;
ROM1[6411]<=26'd1949243; ROM2[6411]<=26'd11124147; ROM3[6411]<=26'd9732225; ROM4[6411]<=26'd23447747;
ROM1[6412]<=26'd1944262; ROM2[6412]<=26'd11124412; ROM3[6412]<=26'd9733210; ROM4[6412]<=26'd23448155;
ROM1[6413]<=26'd1950458; ROM2[6413]<=26'd11127498; ROM3[6413]<=26'd9733935; ROM4[6413]<=26'd23449720;
ROM1[6414]<=26'd1958575; ROM2[6414]<=26'd11127370; ROM3[6414]<=26'd9727945; ROM4[6414]<=26'd23448067;
ROM1[6415]<=26'd1969168; ROM2[6415]<=26'd11126504; ROM3[6415]<=26'd9720436; ROM4[6415]<=26'd23446464;
ROM1[6416]<=26'd1969137; ROM2[6416]<=26'd11124931; ROM3[6416]<=26'd9717762; ROM4[6416]<=26'd23445271;
ROM1[6417]<=26'd1963202; ROM2[6417]<=26'd11125206; ROM3[6417]<=26'd9721827; ROM4[6417]<=26'd23446031;
ROM1[6418]<=26'd1966320; ROM2[6418]<=26'd11132704; ROM3[6418]<=26'd9734595; ROM4[6418]<=26'd23455939;
ROM1[6419]<=26'd1967731; ROM2[6419]<=26'd11136641; ROM3[6419]<=26'd9744249; ROM4[6419]<=26'd23461030;
ROM1[6420]<=26'd1959226; ROM2[6420]<=26'd11132457; ROM3[6420]<=26'd9741978; ROM4[6420]<=26'd23458688;
ROM1[6421]<=26'd1954505; ROM2[6421]<=26'd11126850; ROM3[6421]<=26'd9737418; ROM4[6421]<=26'd23455910;
ROM1[6422]<=26'd1959600; ROM2[6422]<=26'd11125734; ROM3[6422]<=26'd9734590; ROM4[6422]<=26'd23453978;
ROM1[6423]<=26'd1974930; ROM2[6423]<=26'd11129873; ROM3[6423]<=26'd9729365; ROM4[6423]<=26'd23456296;
ROM1[6424]<=26'd1982742; ROM2[6424]<=26'd11130968; ROM3[6424]<=26'd9725769; ROM4[6424]<=26'd23454768;
ROM1[6425]<=26'd1978908; ROM2[6425]<=26'd11131424; ROM3[6425]<=26'd9727903; ROM4[6425]<=26'd23454874;
ROM1[6426]<=26'd1969744; ROM2[6426]<=26'd11131302; ROM3[6426]<=26'd9731777; ROM4[6426]<=26'd23456236;
ROM1[6427]<=26'd1959593; ROM2[6427]<=26'd11128825; ROM3[6427]<=26'd9735225; ROM4[6427]<=26'd23455099;
ROM1[6428]<=26'd1959100; ROM2[6428]<=26'd11135960; ROM3[6428]<=26'd9744601; ROM4[6428]<=26'd23462754;
ROM1[6429]<=26'd1954413; ROM2[6429]<=26'd11134792; ROM3[6429]<=26'd9744674; ROM4[6429]<=26'd23461040;
ROM1[6430]<=26'd1950323; ROM2[6430]<=26'd11127112; ROM3[6430]<=26'd9733520; ROM4[6430]<=26'd23450545;
ROM1[6431]<=26'd1964234; ROM2[6431]<=26'd11129541; ROM3[6431]<=26'd9727812; ROM4[6431]<=26'd23449515;
ROM1[6432]<=26'd1974000; ROM2[6432]<=26'd11127753; ROM3[6432]<=26'd9722633; ROM4[6432]<=26'd23448459;
ROM1[6433]<=26'd1969860; ROM2[6433]<=26'd11126366; ROM3[6433]<=26'd9721139; ROM4[6433]<=26'd23447581;
ROM1[6434]<=26'd1966749; ROM2[6434]<=26'd11129643; ROM3[6434]<=26'd9728057; ROM4[6434]<=26'd23453707;
ROM1[6435]<=26'd1961656; ROM2[6435]<=26'd11128513; ROM3[6435]<=26'd9733325; ROM4[6435]<=26'd23456845;
ROM1[6436]<=26'd1955347; ROM2[6436]<=26'd11127037; ROM3[6436]<=26'd9734361; ROM4[6436]<=26'd23454141;
ROM1[6437]<=26'd1949837; ROM2[6437]<=26'd11127780; ROM3[6437]<=26'd9736886; ROM4[6437]<=26'd23453651;
ROM1[6438]<=26'd1952172; ROM2[6438]<=26'd11127956; ROM3[6438]<=26'd9736418; ROM4[6438]<=26'd23454520;
ROM1[6439]<=26'd1962591; ROM2[6439]<=26'd11129278; ROM3[6439]<=26'd9732726; ROM4[6439]<=26'd23455035;
ROM1[6440]<=26'd1972071; ROM2[6440]<=26'd11128050; ROM3[6440]<=26'd9727567; ROM4[6440]<=26'd23453439;
ROM1[6441]<=26'd1971391; ROM2[6441]<=26'd11125131; ROM3[6441]<=26'd9725032; ROM4[6441]<=26'd23452784;
ROM1[6442]<=26'd1966985; ROM2[6442]<=26'd11125417; ROM3[6442]<=26'd9730387; ROM4[6442]<=26'd23455406;
ROM1[6443]<=26'd1959925; ROM2[6443]<=26'd11123820; ROM3[6443]<=26'd9736427; ROM4[6443]<=26'd23456733;
ROM1[6444]<=26'd1963547; ROM2[6444]<=26'd11130674; ROM3[6444]<=26'd9746500; ROM4[6444]<=26'd23465887;
ROM1[6445]<=26'd1961968; ROM2[6445]<=26'd11133757; ROM3[6445]<=26'd9750359; ROM4[6445]<=26'd23468547;
ROM1[6446]<=26'd1952720; ROM2[6446]<=26'd11126452; ROM3[6446]<=26'd9743768; ROM4[6446]<=26'd23459986;
ROM1[6447]<=26'd1950327; ROM2[6447]<=26'd11119157; ROM3[6447]<=26'd9733707; ROM4[6447]<=26'd23451890;
ROM1[6448]<=26'd1956686; ROM2[6448]<=26'd11115400; ROM3[6448]<=26'd9723700; ROM4[6448]<=26'd23446571;
ROM1[6449]<=26'd1970826; ROM2[6449]<=26'd11123173; ROM3[6449]<=26'd9728006; ROM4[6449]<=26'd23453712;
ROM1[6450]<=26'd1971734; ROM2[6450]<=26'd11125089; ROM3[6450]<=26'd9732668; ROM4[6450]<=26'd23456995;
ROM1[6451]<=26'd1964375; ROM2[6451]<=26'd11123175; ROM3[6451]<=26'd9733274; ROM4[6451]<=26'd23455801;
ROM1[6452]<=26'd1960445; ROM2[6452]<=26'd11121930; ROM3[6452]<=26'd9736692; ROM4[6452]<=26'd23456976;
ROM1[6453]<=26'd1958719; ROM2[6453]<=26'd11124983; ROM3[6453]<=26'd9745098; ROM4[6453]<=26'd23461927;
ROM1[6454]<=26'd1957185; ROM2[6454]<=26'd11126154; ROM3[6454]<=26'd9746704; ROM4[6454]<=26'd23463504;
ROM1[6455]<=26'd1959194; ROM2[6455]<=26'd11124281; ROM3[6455]<=26'd9742847; ROM4[6455]<=26'd23461255;
ROM1[6456]<=26'd1973954; ROM2[6456]<=26'd11130386; ROM3[6456]<=26'd9743163; ROM4[6456]<=26'd23463848;
ROM1[6457]<=26'd1985143; ROM2[6457]<=26'd11131527; ROM3[6457]<=26'd9738358; ROM4[6457]<=26'd23464088;
ROM1[6458]<=26'd1979207; ROM2[6458]<=26'd11126470; ROM3[6458]<=26'd9734672; ROM4[6458]<=26'd23460418;
ROM1[6459]<=26'd1973607; ROM2[6459]<=26'd11126584; ROM3[6459]<=26'd9738344; ROM4[6459]<=26'd23460920;
ROM1[6460]<=26'd1967126; ROM2[6460]<=26'd11126920; ROM3[6460]<=26'd9741182; ROM4[6460]<=26'd23461759;
ROM1[6461]<=26'd1954407; ROM2[6461]<=26'd11120794; ROM3[6461]<=26'd9737572; ROM4[6461]<=26'd23455806;
ROM1[6462]<=26'd1949891; ROM2[6462]<=26'd11120202; ROM3[6462]<=26'd9737094; ROM4[6462]<=26'd23455037;
ROM1[6463]<=26'd1954929; ROM2[6463]<=26'd11123819; ROM3[6463]<=26'd9736502; ROM4[6463]<=26'd23455328;
ROM1[6464]<=26'd1960852; ROM2[6464]<=26'd11120209; ROM3[6464]<=26'd9728526; ROM4[6464]<=26'd23449338;
ROM1[6465]<=26'd1969392; ROM2[6465]<=26'd11116993; ROM3[6465]<=26'd9721088; ROM4[6465]<=26'd23446411;
ROM1[6466]<=26'd1974386; ROM2[6466]<=26'd11122143; ROM3[6466]<=26'd9725628; ROM4[6466]<=26'd23451795;
ROM1[6467]<=26'd1973106; ROM2[6467]<=26'd11129019; ROM3[6467]<=26'd9734116; ROM4[6467]<=26'd23458885;
ROM1[6468]<=26'd1967677; ROM2[6468]<=26'd11129722; ROM3[6468]<=26'd9737380; ROM4[6468]<=26'd23460503;
ROM1[6469]<=26'd1959993; ROM2[6469]<=26'd11124095; ROM3[6469]<=26'd9736427; ROM4[6469]<=26'd23457178;
ROM1[6470]<=26'd1952118; ROM2[6470]<=26'd11121435; ROM3[6470]<=26'd9737346; ROM4[6470]<=26'd23456390;
ROM1[6471]<=26'd1951221; ROM2[6471]<=26'd11122247; ROM3[6471]<=26'd9738305; ROM4[6471]<=26'd23457184;
ROM1[6472]<=26'd1955629; ROM2[6472]<=26'd11121558; ROM3[6472]<=26'd9733945; ROM4[6472]<=26'd23455556;
ROM1[6473]<=26'd1971529; ROM2[6473]<=26'd11127833; ROM3[6473]<=26'd9731962; ROM4[6473]<=26'd23457637;
ROM1[6474]<=26'd1982744; ROM2[6474]<=26'd11132178; ROM3[6474]<=26'd9732702; ROM4[6474]<=26'd23460293;
ROM1[6475]<=26'd1975872; ROM2[6475]<=26'd11127682; ROM3[6475]<=26'd9730165; ROM4[6475]<=26'd23457926;
ROM1[6476]<=26'd1965467; ROM2[6476]<=26'd11124702; ROM3[6476]<=26'd9731117; ROM4[6476]<=26'd23455284;
ROM1[6477]<=26'd1964727; ROM2[6477]<=26'd11129141; ROM3[6477]<=26'd9736881; ROM4[6477]<=26'd23459624;
ROM1[6478]<=26'd1965601; ROM2[6478]<=26'd11134879; ROM3[6478]<=26'd9742234; ROM4[6478]<=26'd23464292;
ROM1[6479]<=26'd1961110; ROM2[6479]<=26'd11132237; ROM3[6479]<=26'd9742556; ROM4[6479]<=26'd23461334;
ROM1[6480]<=26'd1962176; ROM2[6480]<=26'd11128827; ROM3[6480]<=26'd9738408; ROM4[6480]<=26'd23458904;
ROM1[6481]<=26'd1974938; ROM2[6481]<=26'd11130755; ROM3[6481]<=26'd9735324; ROM4[6481]<=26'd23460472;
ROM1[6482]<=26'd1987457; ROM2[6482]<=26'd11134865; ROM3[6482]<=26'd9734187; ROM4[6482]<=26'd23462474;
ROM1[6483]<=26'd1986502; ROM2[6483]<=26'd11138236; ROM3[6483]<=26'd9735671; ROM4[6483]<=26'd23463851;
ROM1[6484]<=26'd1973394; ROM2[6484]<=26'd11132527; ROM3[6484]<=26'd9731117; ROM4[6484]<=26'd23458309;
ROM1[6485]<=26'd1960732; ROM2[6485]<=26'd11124784; ROM3[6485]<=26'd9726648; ROM4[6485]<=26'd23451861;
ROM1[6486]<=26'd1951786; ROM2[6486]<=26'd11119172; ROM3[6486]<=26'd9725253; ROM4[6486]<=26'd23447963;
ROM1[6487]<=26'd1946288; ROM2[6487]<=26'd11117961; ROM3[6487]<=26'd9728032; ROM4[6487]<=26'd23448289;
ROM1[6488]<=26'd1956297; ROM2[6488]<=26'd11126754; ROM3[6488]<=26'd9735859; ROM4[6488]<=26'd23456186;
ROM1[6489]<=26'd1969408; ROM2[6489]<=26'd11130880; ROM3[6489]<=26'd9736887; ROM4[6489]<=26'd23458170;
ROM1[6490]<=26'd1976324; ROM2[6490]<=26'd11127627; ROM3[6490]<=26'd9730066; ROM4[6490]<=26'd23456184;
ROM1[6491]<=26'd1976944; ROM2[6491]<=26'd11128310; ROM3[6491]<=26'd9730152; ROM4[6491]<=26'd23458868;
ROM1[6492]<=26'd1970651; ROM2[6492]<=26'd11126230; ROM3[6492]<=26'd9734000; ROM4[6492]<=26'd23458700;
ROM1[6493]<=26'd1964448; ROM2[6493]<=26'd11127924; ROM3[6493]<=26'd9741136; ROM4[6493]<=26'd23463067;
ROM1[6494]<=26'd1959033; ROM2[6494]<=26'd11129848; ROM3[6494]<=26'd9742537; ROM4[6494]<=26'd23463866;
ROM1[6495]<=26'd1950231; ROM2[6495]<=26'd11123954; ROM3[6495]<=26'd9737299; ROM4[6495]<=26'd23456859;
ROM1[6496]<=26'd1945528; ROM2[6496]<=26'd11119234; ROM3[6496]<=26'd9733365; ROM4[6496]<=26'd23453357;
ROM1[6497]<=26'd1947931; ROM2[6497]<=26'd11115201; ROM3[6497]<=26'd9725965; ROM4[6497]<=26'd23449847;
ROM1[6498]<=26'd1963218; ROM2[6498]<=26'd11118088; ROM3[6498]<=26'd9723406; ROM4[6498]<=26'd23452034;
ROM1[6499]<=26'd1974703; ROM2[6499]<=26'd11123818; ROM3[6499]<=26'd9726903; ROM4[6499]<=26'd23457305;
ROM1[6500]<=26'd1971154; ROM2[6500]<=26'd11124924; ROM3[6500]<=26'd9729704; ROM4[6500]<=26'd23458071;
ROM1[6501]<=26'd1963693; ROM2[6501]<=26'd11125235; ROM3[6501]<=26'd9732848; ROM4[6501]<=26'd23458315;
ROM1[6502]<=26'd1965388; ROM2[6502]<=26'd11133821; ROM3[6502]<=26'd9744798; ROM4[6502]<=26'd23466929;
ROM1[6503]<=26'd1960902; ROM2[6503]<=26'd11133299; ROM3[6503]<=26'd9748860; ROM4[6503]<=26'd23468352;
ROM1[6504]<=26'd1949603; ROM2[6504]<=26'd11124372; ROM3[6504]<=26'd9739393; ROM4[6504]<=26'd23459152;
ROM1[6505]<=26'd1950399; ROM2[6505]<=26'd11122945; ROM3[6505]<=26'd9732341; ROM4[6505]<=26'd23452974;
ROM1[6506]<=26'd1961043; ROM2[6506]<=26'd11123186; ROM3[6506]<=26'd9724671; ROM4[6506]<=26'd23449685;
ROM1[6507]<=26'd1970355; ROM2[6507]<=26'd11124691; ROM3[6507]<=26'd9719149; ROM4[6507]<=26'd23447893;
ROM1[6508]<=26'd1970707; ROM2[6508]<=26'd11128203; ROM3[6508]<=26'd9724596; ROM4[6508]<=26'd23452538;
ROM1[6509]<=26'd1964819; ROM2[6509]<=26'd11128926; ROM3[6509]<=26'd9731514; ROM4[6509]<=26'd23455928;
ROM1[6510]<=26'd1952684; ROM2[6510]<=26'd11121417; ROM3[6510]<=26'd9730739; ROM4[6510]<=26'd23450510;
ROM1[6511]<=26'd1945345; ROM2[6511]<=26'd11117301; ROM3[6511]<=26'd9731157; ROM4[6511]<=26'd23447666;
ROM1[6512]<=26'd1944778; ROM2[6512]<=26'd11119854; ROM3[6512]<=26'd9736069; ROM4[6512]<=26'd23451299;
ROM1[6513]<=26'd1946498; ROM2[6513]<=26'd11119487; ROM3[6513]<=26'd9736696; ROM4[6513]<=26'd23452499;
ROM1[6514]<=26'd1956029; ROM2[6514]<=26'd11120534; ROM3[6514]<=26'd9734919; ROM4[6514]<=26'd23453530;
ROM1[6515]<=26'd1969267; ROM2[6515]<=26'd11123075; ROM3[6515]<=26'd9730827; ROM4[6515]<=26'd23455858;
ROM1[6516]<=26'd1973409; ROM2[6516]<=26'd11125399; ROM3[6516]<=26'd9731164; ROM4[6516]<=26'd23456776;
ROM1[6517]<=26'd1970936; ROM2[6517]<=26'd11128427; ROM3[6517]<=26'd9735458; ROM4[6517]<=26'd23459475;
ROM1[6518]<=26'd1965731; ROM2[6518]<=26'd11128786; ROM3[6518]<=26'd9739677; ROM4[6518]<=26'd23460662;
ROM1[6519]<=26'd1959106; ROM2[6519]<=26'd11127245; ROM3[6519]<=26'd9741525; ROM4[6519]<=26'd23460332;
ROM1[6520]<=26'd1952711; ROM2[6520]<=26'd11125318; ROM3[6520]<=26'd9742742; ROM4[6520]<=26'd23458566;
ROM1[6521]<=26'd1952304; ROM2[6521]<=26'd11124746; ROM3[6521]<=26'd9740717; ROM4[6521]<=26'd23457146;
ROM1[6522]<=26'd1957151; ROM2[6522]<=26'd11124430; ROM3[6522]<=26'd9735877; ROM4[6522]<=26'd23456273;
ROM1[6523]<=26'd1973151; ROM2[6523]<=26'd11128042; ROM3[6523]<=26'd9736144; ROM4[6523]<=26'd23460302;
ROM1[6524]<=26'd1983792; ROM2[6524]<=26'd11132978; ROM3[6524]<=26'd9739338; ROM4[6524]<=26'd23466176;
ROM1[6525]<=26'd1980552; ROM2[6525]<=26'd11134704; ROM3[6525]<=26'd9745022; ROM4[6525]<=26'd23470379;
ROM1[6526]<=26'd1969213; ROM2[6526]<=26'd11130466; ROM3[6526]<=26'd9745904; ROM4[6526]<=26'd23468253;
ROM1[6527]<=26'd1957878; ROM2[6527]<=26'd11123529; ROM3[6527]<=26'd9742712; ROM4[6527]<=26'd23461019;
ROM1[6528]<=26'd1954498; ROM2[6528]<=26'd11127277; ROM3[6528]<=26'd9748705; ROM4[6528]<=26'd23465083;
ROM1[6529]<=26'd1951072; ROM2[6529]<=26'd11128565; ROM3[6529]<=26'd9750073; ROM4[6529]<=26'd23465059;
ROM1[6530]<=26'd1956712; ROM2[6530]<=26'd11128526; ROM3[6530]<=26'd9749940; ROM4[6530]<=26'd23463939;
ROM1[6531]<=26'd1973526; ROM2[6531]<=26'd11132714; ROM3[6531]<=26'd9750086; ROM4[6531]<=26'd23468677;
ROM1[6532]<=26'd1980408; ROM2[6532]<=26'd11128803; ROM3[6532]<=26'd9743320; ROM4[6532]<=26'd23465299;
ROM1[6533]<=26'd1977635; ROM2[6533]<=26'd11125577; ROM3[6533]<=26'd9743348; ROM4[6533]<=26'd23463595;
ROM1[6534]<=26'd1976716; ROM2[6534]<=26'd11130706; ROM3[6534]<=26'd9751105; ROM4[6534]<=26'd23468976;
ROM1[6535]<=26'd1970120; ROM2[6535]<=26'd11130201; ROM3[6535]<=26'd9755471; ROM4[6535]<=26'd23470130;
ROM1[6536]<=26'd1958177; ROM2[6536]<=26'd11122514; ROM3[6536]<=26'd9750508; ROM4[6536]<=26'd23465501;
ROM1[6537]<=26'd1950867; ROM2[6537]<=26'd11119570; ROM3[6537]<=26'd9749385; ROM4[6537]<=26'd23463440;
ROM1[6538]<=26'd1951332; ROM2[6538]<=26'd11119845; ROM3[6538]<=26'd9747715; ROM4[6538]<=26'd23462563;
ROM1[6539]<=26'd1956316; ROM2[6539]<=26'd11117443; ROM3[6539]<=26'd9737421; ROM4[6539]<=26'd23456736;
ROM1[6540]<=26'd1970237; ROM2[6540]<=26'd11119928; ROM3[6540]<=26'd9734613; ROM4[6540]<=26'd23457728;
ROM1[6541]<=26'd1979007; ROM2[6541]<=26'd11126201; ROM3[6541]<=26'd9739336; ROM4[6541]<=26'd23463350;
ROM1[6542]<=26'd1975188; ROM2[6542]<=26'd11128348; ROM3[6542]<=26'd9743677; ROM4[6542]<=26'd23466600;
ROM1[6543]<=26'd1964608; ROM2[6543]<=26'd11124724; ROM3[6543]<=26'd9744259; ROM4[6543]<=26'd23464725;
ROM1[6544]<=26'd1953566; ROM2[6544]<=26'd11119220; ROM3[6544]<=26'd9741101; ROM4[6544]<=26'd23458557;
ROM1[6545]<=26'd1941753; ROM2[6545]<=26'd11111318; ROM3[6545]<=26'd9737666; ROM4[6545]<=26'd23453352;
ROM1[6546]<=26'd1937551; ROM2[6546]<=26'd11105939; ROM3[6546]<=26'd9733281; ROM4[6546]<=26'd23449184;
ROM1[6547]<=26'd1948109; ROM2[6547]<=26'd11111697; ROM3[6547]<=26'd9736543; ROM4[6547]<=26'd23452163;
ROM1[6548]<=26'd1972698; ROM2[6548]<=26'd11124623; ROM3[6548]<=26'd9743082; ROM4[6548]<=26'd23463449;
ROM1[6549]<=26'd1979767; ROM2[6549]<=26'd11127492; ROM3[6549]<=26'd9741373; ROM4[6549]<=26'd23465638;
ROM1[6550]<=26'd1964504; ROM2[6550]<=26'd11118289; ROM3[6550]<=26'd9735565; ROM4[6550]<=26'd23457831;
ROM1[6551]<=26'd1953516; ROM2[6551]<=26'd11115488; ROM3[6551]<=26'd9736616; ROM4[6551]<=26'd23456241;
ROM1[6552]<=26'd1944361; ROM2[6552]<=26'd11113109; ROM3[6552]<=26'd9736341; ROM4[6552]<=26'd23452887;
ROM1[6553]<=26'd1938279; ROM2[6553]<=26'd11110180; ROM3[6553]<=26'd9738653; ROM4[6553]<=26'd23450438;
ROM1[6554]<=26'd1942769; ROM2[6554]<=26'd11117434; ROM3[6554]<=26'd9744985; ROM4[6554]<=26'd23456694;
ROM1[6555]<=26'd1950834; ROM2[6555]<=26'd11120558; ROM3[6555]<=26'd9743668; ROM4[6555]<=26'd23460934;
ROM1[6556]<=26'd1960458; ROM2[6556]<=26'd11118377; ROM3[6556]<=26'd9737726; ROM4[6556]<=26'd23459024;
ROM1[6557]<=26'd1972387; ROM2[6557]<=26'd11122422; ROM3[6557]<=26'd9734684; ROM4[6557]<=26'd23460328;
ROM1[6558]<=26'd1972814; ROM2[6558]<=26'd11124637; ROM3[6558]<=26'd9736352; ROM4[6558]<=26'd23461759;
ROM1[6559]<=26'd1969462; ROM2[6559]<=26'd11128919; ROM3[6559]<=26'd9743518; ROM4[6559]<=26'd23466546;
ROM1[6560]<=26'd1965722; ROM2[6560]<=26'd11131068; ROM3[6560]<=26'd9748183; ROM4[6560]<=26'd23470093;
ROM1[6561]<=26'd1956851; ROM2[6561]<=26'd11125408; ROM3[6561]<=26'd9747193; ROM4[6561]<=26'd23467555;
ROM1[6562]<=26'd1951590; ROM2[6562]<=26'd11122402; ROM3[6562]<=26'd9748596; ROM4[6562]<=26'd23466797;
ROM1[6563]<=26'd1953673; ROM2[6563]<=26'd11122396; ROM3[6563]<=26'd9747816; ROM4[6563]<=26'd23464440;
ROM1[6564]<=26'd1960717; ROM2[6564]<=26'd11122011; ROM3[6564]<=26'd9741962; ROM4[6564]<=26'd23460367;
ROM1[6565]<=26'd1972294; ROM2[6565]<=26'd11124838; ROM3[6565]<=26'd9737463; ROM4[6565]<=26'd23460794;
ROM1[6566]<=26'd1975037; ROM2[6566]<=26'd11125627; ROM3[6566]<=26'd9738390; ROM4[6566]<=26'd23462167;
ROM1[6567]<=26'd1975167; ROM2[6567]<=26'd11129977; ROM3[6567]<=26'd9745213; ROM4[6567]<=26'd23467181;
ROM1[6568]<=26'd1971848; ROM2[6568]<=26'd11132711; ROM3[6568]<=26'd9750771; ROM4[6568]<=26'd23471443;
ROM1[6569]<=26'd1961086; ROM2[6569]<=26'd11128136; ROM3[6569]<=26'd9749796; ROM4[6569]<=26'd23465685;
ROM1[6570]<=26'd1949448; ROM2[6570]<=26'd11123156; ROM3[6570]<=26'd9748494; ROM4[6570]<=26'd23460508;
ROM1[6571]<=26'd1950306; ROM2[6571]<=26'd11125099; ROM3[6571]<=26'd9752050; ROM4[6571]<=26'd23464083;
ROM1[6572]<=26'd1962458; ROM2[6572]<=26'd11130669; ROM3[6572]<=26'd9753450; ROM4[6572]<=26'd23467096;
ROM1[6573]<=26'd1969194; ROM2[6573]<=26'd11125845; ROM3[6573]<=26'd9742699; ROM4[6573]<=26'd23461418;
ROM1[6574]<=26'd1972666; ROM2[6574]<=26'd11124910; ROM3[6574]<=26'd9737821; ROM4[6574]<=26'd23459887;
ROM1[6575]<=26'd1962977; ROM2[6575]<=26'd11119426; ROM3[6575]<=26'd9733962; ROM4[6575]<=26'd23453775;
ROM1[6576]<=26'd1952463; ROM2[6576]<=26'd11116099; ROM3[6576]<=26'd9735354; ROM4[6576]<=26'd23451601;
ROM1[6577]<=26'd1952585; ROM2[6577]<=26'd11121442; ROM3[6577]<=26'd9744581; ROM4[6577]<=26'd23459598;
ROM1[6578]<=26'd1948446; ROM2[6578]<=26'd11122425; ROM3[6578]<=26'd9746776; ROM4[6578]<=26'd23460218;
ROM1[6579]<=26'd1942422; ROM2[6579]<=26'd11119935; ROM3[6579]<=26'd9744170; ROM4[6579]<=26'd23456489;
ROM1[6580]<=26'd1941799; ROM2[6580]<=26'd11115841; ROM3[6580]<=26'd9738109; ROM4[6580]<=26'd23452279;
ROM1[6581]<=26'd1955654; ROM2[6581]<=26'd11119185; ROM3[6581]<=26'd9732465; ROM4[6581]<=26'd23451400;
ROM1[6582]<=26'd1969786; ROM2[6582]<=26'd11124632; ROM3[6582]<=26'd9731449; ROM4[6582]<=26'd23452013;
ROM1[6583]<=26'd1968693; ROM2[6583]<=26'd11125169; ROM3[6583]<=26'd9734128; ROM4[6583]<=26'd23453144;
ROM1[6584]<=26'd1962491; ROM2[6584]<=26'd11125828; ROM3[6584]<=26'd9739144; ROM4[6584]<=26'd23455061;
ROM1[6585]<=26'd1961928; ROM2[6585]<=26'd11129851; ROM3[6585]<=26'd9748410; ROM4[6585]<=26'd23461715;
ROM1[6586]<=26'd1953785; ROM2[6586]<=26'd11124980; ROM3[6586]<=26'd9747511; ROM4[6586]<=26'd23461218;
ROM1[6587]<=26'd1943519; ROM2[6587]<=26'd11117726; ROM3[6587]<=26'd9741671; ROM4[6587]<=26'd23454725;
ROM1[6588]<=26'd1946318; ROM2[6588]<=26'd11118929; ROM3[6588]<=26'd9740585; ROM4[6588]<=26'd23454846;
ROM1[6589]<=26'd1952588; ROM2[6589]<=26'd11117362; ROM3[6589]<=26'd9733307; ROM4[6589]<=26'd23451116;
ROM1[6590]<=26'd1966231; ROM2[6590]<=26'd11120507; ROM3[6590]<=26'd9730262; ROM4[6590]<=26'd23452897;
ROM1[6591]<=26'd1968861; ROM2[6591]<=26'd11123197; ROM3[6591]<=26'd9731884; ROM4[6591]<=26'd23455715;
ROM1[6592]<=26'd1957313; ROM2[6592]<=26'd11116940; ROM3[6592]<=26'd9729015; ROM4[6592]<=26'd23451245;
ROM1[6593]<=26'd1947374; ROM2[6593]<=26'd11112178; ROM3[6593]<=26'd9729109; ROM4[6593]<=26'd23447221;
ROM1[6594]<=26'd1939509; ROM2[6594]<=26'd11110316; ROM3[6594]<=26'd9729051; ROM4[6594]<=26'd23444942;
ROM1[6595]<=26'd1935228; ROM2[6595]<=26'd11110312; ROM3[6595]<=26'd9731554; ROM4[6595]<=26'd23445692;
ROM1[6596]<=26'd1943492; ROM2[6596]<=26'd11117159; ROM3[6596]<=26'd9740679; ROM4[6596]<=26'd23454283;
ROM1[6597]<=26'd1959886; ROM2[6597]<=26'd11128003; ROM3[6597]<=26'd9748528; ROM4[6597]<=26'd23463726;
ROM1[6598]<=26'd1972182; ROM2[6598]<=26'd11127773; ROM3[6598]<=26'd9743021; ROM4[6598]<=26'd23461472;
ROM1[6599]<=26'd1969780; ROM2[6599]<=26'd11120543; ROM3[6599]<=26'd9733899; ROM4[6599]<=26'd23453934;
ROM1[6600]<=26'd1958385; ROM2[6600]<=26'd11115175; ROM3[6600]<=26'd9731076; ROM4[6600]<=26'd23448101;
ROM1[6601]<=26'd1948458; ROM2[6601]<=26'd11111601; ROM3[6601]<=26'd9731728; ROM4[6601]<=26'd23445429;
ROM1[6602]<=26'd1951447; ROM2[6602]<=26'd11118768; ROM3[6602]<=26'd9742013; ROM4[6602]<=26'd23453837;
ROM1[6603]<=26'd1958732; ROM2[6603]<=26'd11131177; ROM3[6603]<=26'd9755608; ROM4[6603]<=26'd23466394;
ROM1[6604]<=26'd1957766; ROM2[6604]<=26'd11131726; ROM3[6604]<=26'd9753259; ROM4[6604]<=26'd23464278;
ROM1[6605]<=26'd1954647; ROM2[6605]<=26'd11123685; ROM3[6605]<=26'd9742603; ROM4[6605]<=26'd23454555;
ROM1[6606]<=26'd1963431; ROM2[6606]<=26'd11122028; ROM3[6606]<=26'd9736520; ROM4[6606]<=26'd23453939;
ROM1[6607]<=26'd1971817; ROM2[6607]<=26'd11120452; ROM3[6607]<=26'd9731793; ROM4[6607]<=26'd23451822;
ROM1[6608]<=26'd1969030; ROM2[6608]<=26'd11119736; ROM3[6608]<=26'd9734951; ROM4[6608]<=26'd23452293;
ROM1[6609]<=26'd1964242; ROM2[6609]<=26'd11121521; ROM3[6609]<=26'd9742020; ROM4[6609]<=26'd23458179;
ROM1[6610]<=26'd1958460; ROM2[6610]<=26'd11121613; ROM3[6610]<=26'd9748179; ROM4[6610]<=26'd23459190;
ROM1[6611]<=26'd1952285; ROM2[6611]<=26'd11120610; ROM3[6611]<=26'd9750604; ROM4[6611]<=26'd23458693;
ROM1[6612]<=26'd1947439; ROM2[6612]<=26'd11119512; ROM3[6612]<=26'd9751608; ROM4[6612]<=26'd23458910;
ROM1[6613]<=26'd1950900; ROM2[6613]<=26'd11121721; ROM3[6613]<=26'd9752476; ROM4[6613]<=26'd23460030;
ROM1[6614]<=26'd1963221; ROM2[6614]<=26'd11126013; ROM3[6614]<=26'd9751119; ROM4[6614]<=26'd23462072;
ROM1[6615]<=26'd1975805; ROM2[6615]<=26'd11127665; ROM3[6615]<=26'd9747363; ROM4[6615]<=26'd23463513;
ROM1[6616]<=26'd1975442; ROM2[6616]<=26'd11124956; ROM3[6616]<=26'd9745775; ROM4[6616]<=26'd23462076;
ROM1[6617]<=26'd1969645; ROM2[6617]<=26'd11124950; ROM3[6617]<=26'd9749927; ROM4[6617]<=26'd23463286;
ROM1[6618]<=26'd1961008; ROM2[6618]<=26'd11123942; ROM3[6618]<=26'd9752338; ROM4[6618]<=26'd23463404;
ROM1[6619]<=26'd1963318; ROM2[6619]<=26'd11131001; ROM3[6619]<=26'd9758835; ROM4[6619]<=26'd23468401;
ROM1[6620]<=26'd1962001; ROM2[6620]<=26'd11133228; ROM3[6620]<=26'd9760802; ROM4[6620]<=26'd23469240;
ROM1[6621]<=26'd1955505; ROM2[6621]<=26'd11127817; ROM3[6621]<=26'd9752732; ROM4[6621]<=26'd23460320;
ROM1[6622]<=26'd1956698; ROM2[6622]<=26'd11123884; ROM3[6622]<=26'd9743286; ROM4[6622]<=26'd23453689;
ROM1[6623]<=26'd1969937; ROM2[6623]<=26'd11124669; ROM3[6623]<=26'd9737839; ROM4[6623]<=26'd23453377;
ROM1[6624]<=26'd1981595; ROM2[6624]<=26'd11131880; ROM3[6624]<=26'd9742696; ROM4[6624]<=26'd23460624;
ROM1[6625]<=26'd1984311; ROM2[6625]<=26'd11139723; ROM3[6625]<=26'd9751990; ROM4[6625]<=26'd23470347;
ROM1[6626]<=26'd1977372; ROM2[6626]<=26'd11136723; ROM3[6626]<=26'd9753270; ROM4[6626]<=26'd23467539;
ROM1[6627]<=26'd1964998; ROM2[6627]<=26'd11128234; ROM3[6627]<=26'd9749712; ROM4[6627]<=26'd23461589;
ROM1[6628]<=26'd1957545; ROM2[6628]<=26'd11129034; ROM3[6628]<=26'd9751917; ROM4[6628]<=26'd23462155;
ROM1[6629]<=26'd1950129; ROM2[6629]<=26'd11123804; ROM3[6629]<=26'd9748564; ROM4[6629]<=26'd23456978;
ROM1[6630]<=26'd1954368; ROM2[6630]<=26'd11121978; ROM3[6630]<=26'd9745657; ROM4[6630]<=26'd23456874;
ROM1[6631]<=26'd1968115; ROM2[6631]<=26'd11125071; ROM3[6631]<=26'd9743952; ROM4[6631]<=26'd23458995;
ROM1[6632]<=26'd1976394; ROM2[6632]<=26'd11123592; ROM3[6632]<=26'd9738678; ROM4[6632]<=26'd23456870;
ROM1[6633]<=26'd1975076; ROM2[6633]<=26'd11122637; ROM3[6633]<=26'd9739829; ROM4[6633]<=26'd23457590;
ROM1[6634]<=26'd1966068; ROM2[6634]<=26'd11122060; ROM3[6634]<=26'd9744432; ROM4[6634]<=26'd23459968;
ROM1[6635]<=26'd1958736; ROM2[6635]<=26'd11121482; ROM3[6635]<=26'd9748836; ROM4[6635]<=26'd23460259;
ROM1[6636]<=26'd1954500; ROM2[6636]<=26'd11122192; ROM3[6636]<=26'd9751342; ROM4[6636]<=26'd23460773;
ROM1[6637]<=26'd1947806; ROM2[6637]<=26'd11119757; ROM3[6637]<=26'd9749250; ROM4[6637]<=26'd23457050;
ROM1[6638]<=26'd1953440; ROM2[6638]<=26'd11124064; ROM3[6638]<=26'd9750000; ROM4[6638]<=26'd23457917;
ROM1[6639]<=26'd1966264; ROM2[6639]<=26'd11130411; ROM3[6639]<=26'd9749519; ROM4[6639]<=26'd23462000;
ROM1[6640]<=26'd1973817; ROM2[6640]<=26'd11127709; ROM3[6640]<=26'd9738208; ROM4[6640]<=26'd23456966;
ROM1[6641]<=26'd1976979; ROM2[6641]<=26'd11129718; ROM3[6641]<=26'd9736162; ROM4[6641]<=26'd23456763;
ROM1[6642]<=26'd1970606; ROM2[6642]<=26'd11127296; ROM3[6642]<=26'd9736212; ROM4[6642]<=26'd23453824;
ROM1[6643]<=26'd1954878; ROM2[6643]<=26'd11118296; ROM3[6643]<=26'd9731297; ROM4[6643]<=26'd23445891;
ROM1[6644]<=26'd1950625; ROM2[6644]<=26'd11115694; ROM3[6644]<=26'd9735071; ROM4[6644]<=26'd23446594;
ROM1[6645]<=26'd1949155; ROM2[6645]<=26'd11117047; ROM3[6645]<=26'd9741096; ROM4[6645]<=26'd23450304;
ROM1[6646]<=26'd1952094; ROM2[6646]<=26'd11122279; ROM3[6646]<=26'd9745315; ROM4[6646]<=26'd23454459;
ROM1[6647]<=26'd1967755; ROM2[6647]<=26'd11130796; ROM3[6647]<=26'd9749377; ROM4[6647]<=26'd23461025;
ROM1[6648]<=26'd1979497; ROM2[6648]<=26'd11130752; ROM3[6648]<=26'd9743226; ROM4[6648]<=26'd23460146;
ROM1[6649]<=26'd1985046; ROM2[6649]<=26'd11131031; ROM3[6649]<=26'd9740530; ROM4[6649]<=26'd23461415;
ROM1[6650]<=26'd1978873; ROM2[6650]<=26'd11129088; ROM3[6650]<=26'd9741206; ROM4[6650]<=26'd23460725;
ROM1[6651]<=26'd1964464; ROM2[6651]<=26'd11122109; ROM3[6651]<=26'd9739516; ROM4[6651]<=26'd23455751;
ROM1[6652]<=26'd1960048; ROM2[6652]<=26'd11125768; ROM3[6652]<=26'd9745616; ROM4[6652]<=26'd23459128;
ROM1[6653]<=26'd1954126; ROM2[6653]<=26'd11124847; ROM3[6653]<=26'd9749496; ROM4[6653]<=26'd23459103;
ROM1[6654]<=26'd1952213; ROM2[6654]<=26'd11126211; ROM3[6654]<=26'd9750691; ROM4[6654]<=26'd23459729;
ROM1[6655]<=26'd1958918; ROM2[6655]<=26'd11130256; ROM3[6655]<=26'd9751337; ROM4[6655]<=26'd23462823;
ROM1[6656]<=26'd1970232; ROM2[6656]<=26'd11129917; ROM3[6656]<=26'd9746270; ROM4[6656]<=26'd23460983;
ROM1[6657]<=26'd1978147; ROM2[6657]<=26'd11130701; ROM3[6657]<=26'd9739059; ROM4[6657]<=26'd23458329;
ROM1[6658]<=26'd1973287; ROM2[6658]<=26'd11127884; ROM3[6658]<=26'd9738250; ROM4[6658]<=26'd23456368;
ROM1[6659]<=26'd1966353; ROM2[6659]<=26'd11128282; ROM3[6659]<=26'd9740598; ROM4[6659]<=26'd23456190;
ROM1[6660]<=26'd1959966; ROM2[6660]<=26'd11130129; ROM3[6660]<=26'd9744112; ROM4[6660]<=26'd23457456;
ROM1[6661]<=26'd1956084; ROM2[6661]<=26'd11129482; ROM3[6661]<=26'd9748226; ROM4[6661]<=26'd23458529;
ROM1[6662]<=26'd1954286; ROM2[6662]<=26'd11129737; ROM3[6662]<=26'd9751165; ROM4[6662]<=26'd23460616;
ROM1[6663]<=26'd1959437; ROM2[6663]<=26'd11131476; ROM3[6663]<=26'd9753457; ROM4[6663]<=26'd23463392;
ROM1[6664]<=26'd1968532; ROM2[6664]<=26'd11131410; ROM3[6664]<=26'd9748296; ROM4[6664]<=26'd23461586;
ROM1[6665]<=26'd1975277; ROM2[6665]<=26'd11128798; ROM3[6665]<=26'd9739257; ROM4[6665]<=26'd23456751;
ROM1[6666]<=26'd1975981; ROM2[6666]<=26'd11127467; ROM3[6666]<=26'd9738034; ROM4[6666]<=26'd23454881;
ROM1[6667]<=26'd1972330; ROM2[6667]<=26'd11127466; ROM3[6667]<=26'd9742393; ROM4[6667]<=26'd23456605;
ROM1[6668]<=26'd1967211; ROM2[6668]<=26'd11128167; ROM3[6668]<=26'd9748415; ROM4[6668]<=26'd23459797;
ROM1[6669]<=26'd1965016; ROM2[6669]<=26'd11132733; ROM3[6669]<=26'd9755546; ROM4[6669]<=26'd23466315;
ROM1[6670]<=26'd1953299; ROM2[6670]<=26'd11127733; ROM3[6670]<=26'd9751862; ROM4[6670]<=26'd23461216;
ROM1[6671]<=26'd1946307; ROM2[6671]<=26'd11120158; ROM3[6671]<=26'd9744338; ROM4[6671]<=26'd23450845;
ROM1[6672]<=26'd1953428; ROM2[6672]<=26'd11118760; ROM3[6672]<=26'd9740025; ROM4[6672]<=26'd23448160;
ROM1[6673]<=26'd1966054; ROM2[6673]<=26'd11119032; ROM3[6673]<=26'd9736145; ROM4[6673]<=26'd23448991;
ROM1[6674]<=26'd1971925; ROM2[6674]<=26'd11119488; ROM3[6674]<=26'd9736241; ROM4[6674]<=26'd23450743;
ROM1[6675]<=26'd1965428; ROM2[6675]<=26'd11119611; ROM3[6675]<=26'd9735841; ROM4[6675]<=26'd23451564;
ROM1[6676]<=26'd1960356; ROM2[6676]<=26'd11123530; ROM3[6676]<=26'd9741627; ROM4[6676]<=26'd23454364;
ROM1[6677]<=26'd1958841; ROM2[6677]<=26'd11127100; ROM3[6677]<=26'd9747250; ROM4[6677]<=26'd23455800;
ROM1[6678]<=26'd1950977; ROM2[6678]<=26'd11125704; ROM3[6678]<=26'd9747963; ROM4[6678]<=26'd23454405;
ROM1[6679]<=26'd1947376; ROM2[6679]<=26'd11124611; ROM3[6679]<=26'd9748252; ROM4[6679]<=26'd23452620;
ROM1[6680]<=26'd1957006; ROM2[6680]<=26'd11127843; ROM3[6680]<=26'd9749203; ROM4[6680]<=26'd23455837;
ROM1[6681]<=26'd1966348; ROM2[6681]<=26'd11127255; ROM3[6681]<=26'd9742818; ROM4[6681]<=26'd23453970;
ROM1[6682]<=26'd1970124; ROM2[6682]<=26'd11123592; ROM3[6682]<=26'd9733467; ROM4[6682]<=26'd23449603;
ROM1[6683]<=26'd1967014; ROM2[6683]<=26'd11122630; ROM3[6683]<=26'd9732965; ROM4[6683]<=26'd23448195;
ROM1[6684]<=26'd1958771; ROM2[6684]<=26'd11119821; ROM3[6684]<=26'd9733639; ROM4[6684]<=26'd23446240;
ROM1[6685]<=26'd1953240; ROM2[6685]<=26'd11119292; ROM3[6685]<=26'd9736185; ROM4[6685]<=26'd23446691;
ROM1[6686]<=26'd1950796; ROM2[6686]<=26'd11122865; ROM3[6686]<=26'd9740594; ROM4[6686]<=26'd23450595;
ROM1[6687]<=26'd1944987; ROM2[6687]<=26'd11122713; ROM3[6687]<=26'd9742081; ROM4[6687]<=26'd23450971;
ROM1[6688]<=26'd1942767; ROM2[6688]<=26'd11120968; ROM3[6688]<=26'd9740132; ROM4[6688]<=26'd23449152;
ROM1[6689]<=26'd1950520; ROM2[6689]<=26'd11120620; ROM3[6689]<=26'd9734867; ROM4[6689]<=26'd23447898;
ROM1[6690]<=26'd1965800; ROM2[6690]<=26'd11123442; ROM3[6690]<=26'd9731240; ROM4[6690]<=26'd23448437;
ROM1[6691]<=26'd1968517; ROM2[6691]<=26'd11125382; ROM3[6691]<=26'd9731722; ROM4[6691]<=26'd23450198;
ROM1[6692]<=26'd1960903; ROM2[6692]<=26'd11124602; ROM3[6692]<=26'd9734856; ROM4[6692]<=26'd23451504;
ROM1[6693]<=26'd1954053; ROM2[6693]<=26'd11123412; ROM3[6693]<=26'd9738589; ROM4[6693]<=26'd23451475;
ROM1[6694]<=26'd1951284; ROM2[6694]<=26'd11124300; ROM3[6694]<=26'd9741036; ROM4[6694]<=26'd23452053;
ROM1[6695]<=26'd1944115; ROM2[6695]<=26'd11120058; ROM3[6695]<=26'd9740508; ROM4[6695]<=26'd23449407;
ROM1[6696]<=26'd1940836; ROM2[6696]<=26'd11117169; ROM3[6696]<=26'd9736216; ROM4[6696]<=26'd23445289;
ROM1[6697]<=26'd1946328; ROM2[6697]<=26'd11117516; ROM3[6697]<=26'd9729721; ROM4[6697]<=26'd23441843;
ROM1[6698]<=26'd1957193; ROM2[6698]<=26'd11118454; ROM3[6698]<=26'd9725777; ROM4[6698]<=26'd23441707;
ROM1[6699]<=26'd1966801; ROM2[6699]<=26'd11122404; ROM3[6699]<=26'd9727409; ROM4[6699]<=26'd23445488;
ROM1[6700]<=26'd1967062; ROM2[6700]<=26'd11124987; ROM3[6700]<=26'd9732804; ROM4[6700]<=26'd23449632;
ROM1[6701]<=26'd1959601; ROM2[6701]<=26'd11125147; ROM3[6701]<=26'd9735836; ROM4[6701]<=26'd23449426;
ROM1[6702]<=26'd1956318; ROM2[6702]<=26'd11126455; ROM3[6702]<=26'd9739294; ROM4[6702]<=26'd23449488;
ROM1[6703]<=26'd1949234; ROM2[6703]<=26'd11121816; ROM3[6703]<=26'd9740800; ROM4[6703]<=26'd23448297;
ROM1[6704]<=26'd1937223; ROM2[6704]<=26'd11112106; ROM3[6704]<=26'd9733546; ROM4[6704]<=26'd23440201;
ROM1[6705]<=26'd1941471; ROM2[6705]<=26'd11112661; ROM3[6705]<=26'd9731850; ROM4[6705]<=26'd23439669;
ROM1[6706]<=26'd1955175; ROM2[6706]<=26'd11115318; ROM3[6706]<=26'd9728902; ROM4[6706]<=26'd23441287;
ROM1[6707]<=26'd1966289; ROM2[6707]<=26'd11120512; ROM3[6707]<=26'd9727378; ROM4[6707]<=26'd23444532;
ROM1[6708]<=26'd1967280; ROM2[6708]<=26'd11124600; ROM3[6708]<=26'd9730626; ROM4[6708]<=26'd23446988;
ROM1[6709]<=26'd1958019; ROM2[6709]<=26'd11121380; ROM3[6709]<=26'd9732311; ROM4[6709]<=26'd23446989;
ROM1[6710]<=26'd1953787; ROM2[6710]<=26'd11123139; ROM3[6710]<=26'd9738520; ROM4[6710]<=26'd23450545;
ROM1[6711]<=26'd1953981; ROM2[6711]<=26'd11126605; ROM3[6711]<=26'd9743319; ROM4[6711]<=26'd23453576;
ROM1[6712]<=26'd1950977; ROM2[6712]<=26'd11127746; ROM3[6712]<=26'd9745125; ROM4[6712]<=26'd23454581;
ROM1[6713]<=26'd1955750; ROM2[6713]<=26'd11130979; ROM3[6713]<=26'd9748257; ROM4[6713]<=26'd23458331;
ROM1[6714]<=26'd1965532; ROM2[6714]<=26'd11130769; ROM3[6714]<=26'd9745755; ROM4[6714]<=26'd23458976;
ROM1[6715]<=26'd1974850; ROM2[6715]<=26'd11128153; ROM3[6715]<=26'd9739435; ROM4[6715]<=26'd23457312;
ROM1[6716]<=26'd1977230; ROM2[6716]<=26'd11127626; ROM3[6716]<=26'd9739236; ROM4[6716]<=26'd23458497;
ROM1[6717]<=26'd1973582; ROM2[6717]<=26'd11129863; ROM3[6717]<=26'd9743059; ROM4[6717]<=26'd23460451;
ROM1[6718]<=26'd1968421; ROM2[6718]<=26'd11131316; ROM3[6718]<=26'd9748872; ROM4[6718]<=26'd23462690;
ROM1[6719]<=26'd1964660; ROM2[6719]<=26'd11132199; ROM3[6719]<=26'd9751645; ROM4[6719]<=26'd23463466;
ROM1[6720]<=26'd1955681; ROM2[6720]<=26'd11129712; ROM3[6720]<=26'd9751391; ROM4[6720]<=26'd23461940;
ROM1[6721]<=26'd1953916; ROM2[6721]<=26'd11126877; ROM3[6721]<=26'd9751145; ROM4[6721]<=26'd23460043;
ROM1[6722]<=26'd1964610; ROM2[6722]<=26'd11129948; ROM3[6722]<=26'd9748977; ROM4[6722]<=26'd23461038;
ROM1[6723]<=26'd1977367; ROM2[6723]<=26'd11132020; ROM3[6723]<=26'd9743474; ROM4[6723]<=26'd23462410;
ROM1[6724]<=26'd1986432; ROM2[6724]<=26'd11135573; ROM3[6724]<=26'd9744853; ROM4[6724]<=26'd23463901;
ROM1[6725]<=26'd1991035; ROM2[6725]<=26'd11144868; ROM3[6725]<=26'd9754986; ROM4[6725]<=26'd23471811;
ROM1[6726]<=26'd1982768; ROM2[6726]<=26'd11145231; ROM3[6726]<=26'd9757779; ROM4[6726]<=26'd23472528;
ROM1[6727]<=26'd1965647; ROM2[6727]<=26'd11133915; ROM3[6727]<=26'd9749760; ROM4[6727]<=26'd23461507;
ROM1[6728]<=26'd1954096; ROM2[6728]<=26'd11127249; ROM3[6728]<=26'd9745705; ROM4[6728]<=26'd23456768;
ROM1[6729]<=26'd1949921; ROM2[6729]<=26'd11124851; ROM3[6729]<=26'd9744608; ROM4[6729]<=26'd23455072;
ROM1[6730]<=26'd1952208; ROM2[6730]<=26'd11122427; ROM3[6730]<=26'd9740848; ROM4[6730]<=26'd23453409;
ROM1[6731]<=26'd1966135; ROM2[6731]<=26'd11127475; ROM3[6731]<=26'd9739376; ROM4[6731]<=26'd23456258;
ROM1[6732]<=26'd1976083; ROM2[6732]<=26'd11130692; ROM3[6732]<=26'd9737597; ROM4[6732]<=26'd23458195;
ROM1[6733]<=26'd1967373; ROM2[6733]<=26'd11124475; ROM3[6733]<=26'd9733307; ROM4[6733]<=26'd23453968;
ROM1[6734]<=26'd1959343; ROM2[6734]<=26'd11121619; ROM3[6734]<=26'd9735087; ROM4[6734]<=26'd23451737;
ROM1[6735]<=26'd1958111; ROM2[6735]<=26'd11124119; ROM3[6735]<=26'd9741312; ROM4[6735]<=26'd23454779;
ROM1[6736]<=26'd1960161; ROM2[6736]<=26'd11131214; ROM3[6736]<=26'd9752298; ROM4[6736]<=26'd23464260;
ROM1[6737]<=26'd1957854; ROM2[6737]<=26'd11131719; ROM3[6737]<=26'd9755211; ROM4[6737]<=26'd23467562;
ROM1[6738]<=26'd1956107; ROM2[6738]<=26'd11128056; ROM3[6738]<=26'd9749799; ROM4[6738]<=26'd23462979;
ROM1[6739]<=26'd1964107; ROM2[6739]<=26'd11127806; ROM3[6739]<=26'd9745950; ROM4[6739]<=26'd23462534;
ROM1[6740]<=26'd1975665; ROM2[6740]<=26'd11127209; ROM3[6740]<=26'd9738872; ROM4[6740]<=26'd23459752;
ROM1[6741]<=26'd1977145; ROM2[6741]<=26'd11127067; ROM3[6741]<=26'd9737018; ROM4[6741]<=26'd23458346;
ROM1[6742]<=26'd1971447; ROM2[6742]<=26'd11127676; ROM3[6742]<=26'd9739832; ROM4[6742]<=26'd23459996;
ROM1[6743]<=26'd1966319; ROM2[6743]<=26'd11127660; ROM3[6743]<=26'd9743743; ROM4[6743]<=26'd23460273;
ROM1[6744]<=26'd1965680; ROM2[6744]<=26'd11130845; ROM3[6744]<=26'd9749502; ROM4[6744]<=26'd23463970;
ROM1[6745]<=26'd1969833; ROM2[6745]<=26'd11140642; ROM3[6745]<=26'd9761605; ROM4[6745]<=26'd23473261;
ROM1[6746]<=26'd1972156; ROM2[6746]<=26'd11143166; ROM3[6746]<=26'd9764608; ROM4[6746]<=26'd23476934;
ROM1[6747]<=26'd1972551; ROM2[6747]<=26'd11137441; ROM3[6747]<=26'd9756342; ROM4[6747]<=26'd23471985;
ROM1[6748]<=26'd1978240; ROM2[6748]<=26'd11131453; ROM3[6748]<=26'd9746590; ROM4[6748]<=26'd23464498;
ROM1[6749]<=26'd1974017; ROM2[6749]<=26'd11122499; ROM3[6749]<=26'd9734389; ROM4[6749]<=26'd23454973;
ROM1[6750]<=26'd1966647; ROM2[6750]<=26'd11120300; ROM3[6750]<=26'd9732085; ROM4[6750]<=26'd23452514;
ROM1[6751]<=26'd1964552; ROM2[6751]<=26'd11125975; ROM3[6751]<=26'd9738135; ROM4[6751]<=26'd23458490;
ROM1[6752]<=26'd1961231; ROM2[6752]<=26'd11128313; ROM3[6752]<=26'd9740800; ROM4[6752]<=26'd23460182;
ROM1[6753]<=26'd1953176; ROM2[6753]<=26'd11125632; ROM3[6753]<=26'd9743017; ROM4[6753]<=26'd23457346;
ROM1[6754]<=26'd1949261; ROM2[6754]<=26'd11123663; ROM3[6754]<=26'd9744807; ROM4[6754]<=26'd23456680;
ROM1[6755]<=26'd1953331; ROM2[6755]<=26'd11123526; ROM3[6755]<=26'd9740619; ROM4[6755]<=26'd23454813;
ROM1[6756]<=26'd1959669; ROM2[6756]<=26'd11120357; ROM3[6756]<=26'd9730322; ROM4[6756]<=26'd23448736;
ROM1[6757]<=26'd1967057; ROM2[6757]<=26'd11120082; ROM3[6757]<=26'd9723627; ROM4[6757]<=26'd23447328;
ROM1[6758]<=26'd1966218; ROM2[6758]<=26'd11120310; ROM3[6758]<=26'd9726428; ROM4[6758]<=26'd23449226;
ROM1[6759]<=26'd1960659; ROM2[6759]<=26'd11122582; ROM3[6759]<=26'd9732873; ROM4[6759]<=26'd23450298;
ROM1[6760]<=26'd1956166; ROM2[6760]<=26'd11125159; ROM3[6760]<=26'd9738269; ROM4[6760]<=26'd23452902;
ROM1[6761]<=26'd1951595; ROM2[6761]<=26'd11125912; ROM3[6761]<=26'd9741296; ROM4[6761]<=26'd23454219;
ROM1[6762]<=26'd1949635; ROM2[6762]<=26'd11128457; ROM3[6762]<=26'd9743621; ROM4[6762]<=26'd23456469;
ROM1[6763]<=26'd1952356; ROM2[6763]<=26'd11127977; ROM3[6763]<=26'd9743154; ROM4[6763]<=26'd23457088;
ROM1[6764]<=26'd1963312; ROM2[6764]<=26'd11130151; ROM3[6764]<=26'd9741421; ROM4[6764]<=26'd23459014;
ROM1[6765]<=26'd1979121; ROM2[6765]<=26'd11133868; ROM3[6765]<=26'd9740926; ROM4[6765]<=26'd23463122;
ROM1[6766]<=26'd1979417; ROM2[6766]<=26'd11132532; ROM3[6766]<=26'd9739534; ROM4[6766]<=26'd23460376;
ROM1[6767]<=26'd1974197; ROM2[6767]<=26'd11133802; ROM3[6767]<=26'd9742329; ROM4[6767]<=26'd23462323;
ROM1[6768]<=26'd1965612; ROM2[6768]<=26'd11132415; ROM3[6768]<=26'd9744047; ROM4[6768]<=26'd23460911;
ROM1[6769]<=26'd1956142; ROM2[6769]<=26'd11130262; ROM3[6769]<=26'd9742530; ROM4[6769]<=26'd23458007;
ROM1[6770]<=26'd1951432; ROM2[6770]<=26'd11131548; ROM3[6770]<=26'd9745048; ROM4[6770]<=26'd23460807;
ROM1[6771]<=26'd1953868; ROM2[6771]<=26'd11134638; ROM3[6771]<=26'd9750075; ROM4[6771]<=26'd23462637;
ROM1[6772]<=26'd1963665; ROM2[6772]<=26'd11135886; ROM3[6772]<=26'd9749919; ROM4[6772]<=26'd23463456;
ROM1[6773]<=26'd1973997; ROM2[6773]<=26'd11132877; ROM3[6773]<=26'd9741894; ROM4[6773]<=26'd23460949;
ROM1[6774]<=26'd1973641; ROM2[6774]<=26'd11128527; ROM3[6774]<=26'd9736295; ROM4[6774]<=26'd23457128;
ROM1[6775]<=26'd1968705; ROM2[6775]<=26'd11127407; ROM3[6775]<=26'd9738697; ROM4[6775]<=26'd23458175;
ROM1[6776]<=26'd1965806; ROM2[6776]<=26'd11131503; ROM3[6776]<=26'd9744988; ROM4[6776]<=26'd23464373;
ROM1[6777]<=26'd1961411; ROM2[6777]<=26'd11132099; ROM3[6777]<=26'd9748525; ROM4[6777]<=26'd23464624;
ROM1[6778]<=26'd1953983; ROM2[6778]<=26'd11129787; ROM3[6778]<=26'd9750730; ROM4[6778]<=26'd23463680;
ROM1[6779]<=26'd1948567; ROM2[6779]<=26'd11126380; ROM3[6779]<=26'd9750929; ROM4[6779]<=26'd23464124;
ROM1[6780]<=26'd1950008; ROM2[6780]<=26'd11123594; ROM3[6780]<=26'd9746895; ROM4[6780]<=26'd23461314;
ROM1[6781]<=26'd1964908; ROM2[6781]<=26'd11127737; ROM3[6781]<=26'd9742494; ROM4[6781]<=26'd23463086;
ROM1[6782]<=26'd1976271; ROM2[6782]<=26'd11132174; ROM3[6782]<=26'd9739464; ROM4[6782]<=26'd23465573;
ROM1[6783]<=26'd1972585; ROM2[6783]<=26'd11131766; ROM3[6783]<=26'd9738974; ROM4[6783]<=26'd23465349;
ROM1[6784]<=26'd1965897; ROM2[6784]<=26'd11129821; ROM3[6784]<=26'd9741909; ROM4[6784]<=26'd23466096;
ROM1[6785]<=26'd1961963; ROM2[6785]<=26'd11128967; ROM3[6785]<=26'd9747961; ROM4[6785]<=26'd23469187;
ROM1[6786]<=26'd1960813; ROM2[6786]<=26'd11130127; ROM3[6786]<=26'd9751777; ROM4[6786]<=26'd23470445;
ROM1[6787]<=26'd1956441; ROM2[6787]<=26'd11128632; ROM3[6787]<=26'd9751987; ROM4[6787]<=26'd23468541;
ROM1[6788]<=26'd1955766; ROM2[6788]<=26'd11126863; ROM3[6788]<=26'd9748419; ROM4[6788]<=26'd23467505;
ROM1[6789]<=26'd1970782; ROM2[6789]<=26'd11136453; ROM3[6789]<=26'd9751024; ROM4[6789]<=26'd23473358;
ROM1[6790]<=26'd1998170; ROM2[6790]<=26'd11155143; ROM3[6790]<=26'd9763380; ROM4[6790]<=26'd23489080;
ROM1[6791]<=26'd1996744; ROM2[6791]<=26'd11152126; ROM3[6791]<=26'd9760512; ROM4[6791]<=26'd23485723;
ROM1[6792]<=26'd1978319; ROM2[6792]<=26'd11137267; ROM3[6792]<=26'd9749832; ROM4[6792]<=26'd23472061;
ROM1[6793]<=26'd1964260; ROM2[6793]<=26'd11127163; ROM3[6793]<=26'd9745975; ROM4[6793]<=26'd23464938;
ROM1[6794]<=26'd1951660; ROM2[6794]<=26'd11118775; ROM3[6794]<=26'd9742361; ROM4[6794]<=26'd23457606;
ROM1[6795]<=26'd1945367; ROM2[6795]<=26'd11118970; ROM3[6795]<=26'd9744190; ROM4[6795]<=26'd23455022;
ROM1[6796]<=26'd1949701; ROM2[6796]<=26'd11125870; ROM3[6796]<=26'd9749013; ROM4[6796]<=26'd23458941;
ROM1[6797]<=26'd1958569; ROM2[6797]<=26'd11129543; ROM3[6797]<=26'd9746800; ROM4[6797]<=26'd23459264;
ROM1[6798]<=26'd1967910; ROM2[6798]<=26'd11127297; ROM3[6798]<=26'd9739556; ROM4[6798]<=26'd23456528;
ROM1[6799]<=26'd1976856; ROM2[6799]<=26'd11130259; ROM3[6799]<=26'd9740769; ROM4[6799]<=26'd23461166;
ROM1[6800]<=26'd1975834; ROM2[6800]<=26'd11133823; ROM3[6800]<=26'd9745156; ROM4[6800]<=26'd23464147;
ROM1[6801]<=26'd1962277; ROM2[6801]<=26'd11128341; ROM3[6801]<=26'd9743389; ROM4[6801]<=26'd23458933;
ROM1[6802]<=26'd1954531; ROM2[6802]<=26'd11126120; ROM3[6802]<=26'd9741755; ROM4[6802]<=26'd23457141;
ROM1[6803]<=26'd1950061; ROM2[6803]<=26'd11127579; ROM3[6803]<=26'd9743901; ROM4[6803]<=26'd23457515;
ROM1[6804]<=26'd1947922; ROM2[6804]<=26'd11127905; ROM3[6804]<=26'd9745827; ROM4[6804]<=26'd23457636;
ROM1[6805]<=26'd1952489; ROM2[6805]<=26'd11125850; ROM3[6805]<=26'd9742970; ROM4[6805]<=26'd23456283;
ROM1[6806]<=26'd1961535; ROM2[6806]<=26'd11122701; ROM3[6806]<=26'd9734024; ROM4[6806]<=26'd23451099;
ROM1[6807]<=26'd1969746; ROM2[6807]<=26'd11122794; ROM3[6807]<=26'd9728630; ROM4[6807]<=26'd23450678;
ROM1[6808]<=26'd1970736; ROM2[6808]<=26'd11125806; ROM3[6808]<=26'd9732246; ROM4[6808]<=26'd23453357;
ROM1[6809]<=26'd1968563; ROM2[6809]<=26'd11130126; ROM3[6809]<=26'd9738496; ROM4[6809]<=26'd23457322;
ROM1[6810]<=26'd1959970; ROM2[6810]<=26'd11128928; ROM3[6810]<=26'd9740235; ROM4[6810]<=26'd23457229;
ROM1[6811]<=26'd1951179; ROM2[6811]<=26'd11126243; ROM3[6811]<=26'd9739053; ROM4[6811]<=26'd23454712;
ROM1[6812]<=26'd1949657; ROM2[6812]<=26'd11129092; ROM3[6812]<=26'd9742560; ROM4[6812]<=26'd23456835;
ROM1[6813]<=26'd1951922; ROM2[6813]<=26'd11130651; ROM3[6813]<=26'd9741437; ROM4[6813]<=26'd23457803;
ROM1[6814]<=26'd1960633; ROM2[6814]<=26'd11130177; ROM3[6814]<=26'd9734840; ROM4[6814]<=26'd23453694;
ROM1[6815]<=26'd1974382; ROM2[6815]<=26'd11131715; ROM3[6815]<=26'd9731470; ROM4[6815]<=26'd23454147;
ROM1[6816]<=26'd1975907; ROM2[6816]<=26'd11131354; ROM3[6816]<=26'd9733712; ROM4[6816]<=26'd23456345;
ROM1[6817]<=26'd1970120; ROM2[6817]<=26'd11130692; ROM3[6817]<=26'd9737939; ROM4[6817]<=26'd23457322;
ROM1[6818]<=26'd1963651; ROM2[6818]<=26'd11131138; ROM3[6818]<=26'd9741889; ROM4[6818]<=26'd23458990;
ROM1[6819]<=26'd1958105; ROM2[6819]<=26'd11129273; ROM3[6819]<=26'd9744029; ROM4[6819]<=26'd23458153;
ROM1[6820]<=26'd1953339; ROM2[6820]<=26'd11129029; ROM3[6820]<=26'd9744845; ROM4[6820]<=26'd23458848;
ROM1[6821]<=26'd1964126; ROM2[6821]<=26'd11140035; ROM3[6821]<=26'd9756250; ROM4[6821]<=26'd23468940;
ROM1[6822]<=26'd1975273; ROM2[6822]<=26'd11144125; ROM3[6822]<=26'd9758563; ROM4[6822]<=26'd23472048;
ROM1[6823]<=26'd1978973; ROM2[6823]<=26'd11136726; ROM3[6823]<=26'd9743980; ROM4[6823]<=26'd23465483;
ROM1[6824]<=26'd1987883; ROM2[6824]<=26'd11139877; ROM3[6824]<=26'd9744993; ROM4[6824]<=26'd23469207;
ROM1[6825]<=26'd1975265; ROM2[6825]<=26'd11130823; ROM3[6825]<=26'd9737685; ROM4[6825]<=26'd23460966;
ROM1[6826]<=26'd1959550; ROM2[6826]<=26'd11121220; ROM3[6826]<=26'd9731991; ROM4[6826]<=26'd23453223;
ROM1[6827]<=26'd1958132; ROM2[6827]<=26'd11124912; ROM3[6827]<=26'd9738326; ROM4[6827]<=26'd23457203;
ROM1[6828]<=26'd1947392; ROM2[6828]<=26'd11121712; ROM3[6828]<=26'd9736711; ROM4[6828]<=26'd23453513;
ROM1[6829]<=26'd1941507; ROM2[6829]<=26'd11117996; ROM3[6829]<=26'd9736079; ROM4[6829]<=26'd23450438;
ROM1[6830]<=26'd1948724; ROM2[6830]<=26'd11120031; ROM3[6830]<=26'd9734486; ROM4[6830]<=26'd23451866;
ROM1[6831]<=26'd1962321; ROM2[6831]<=26'd11124968; ROM3[6831]<=26'd9731693; ROM4[6831]<=26'd23452056;
ROM1[6832]<=26'd1968406; ROM2[6832]<=26'd11122142; ROM3[6832]<=26'd9726780; ROM4[6832]<=26'd23448250;
ROM1[6833]<=26'd1964602; ROM2[6833]<=26'd11119970; ROM3[6833]<=26'd9725711; ROM4[6833]<=26'd23447146;
ROM1[6834]<=26'd1961784; ROM2[6834]<=26'd11122949; ROM3[6834]<=26'd9731849; ROM4[6834]<=26'd23449951;
ROM1[6835]<=26'd1961811; ROM2[6835]<=26'd11128296; ROM3[6835]<=26'd9738946; ROM4[6835]<=26'd23455950;
ROM1[6836]<=26'd1960495; ROM2[6836]<=26'd11132327; ROM3[6836]<=26'd9743679; ROM4[6836]<=26'd23461034;
ROM1[6837]<=26'd1958022; ROM2[6837]<=26'd11133768; ROM3[6837]<=26'd9747460; ROM4[6837]<=26'd23462787;
ROM1[6838]<=26'd1962629; ROM2[6838]<=26'd11137132; ROM3[6838]<=26'd9749523; ROM4[6838]<=26'd23465838;
ROM1[6839]<=26'd1974102; ROM2[6839]<=26'd11139053; ROM3[6839]<=26'd9749407; ROM4[6839]<=26'd23468171;
ROM1[6840]<=26'd1983183; ROM2[6840]<=26'd11134939; ROM3[6840]<=26'd9741131; ROM4[6840]<=26'd23463899;
ROM1[6841]<=26'd1981050; ROM2[6841]<=26'd11132880; ROM3[6841]<=26'd9735572; ROM4[6841]<=26'd23460449;
ROM1[6842]<=26'd1972925; ROM2[6842]<=26'd11130875; ROM3[6842]<=26'd9738109; ROM4[6842]<=26'd23460987;
ROM1[6843]<=26'd1964412; ROM2[6843]<=26'd11128164; ROM3[6843]<=26'd9740854; ROM4[6843]<=26'd23459563;
ROM1[6844]<=26'd1960608; ROM2[6844]<=26'd11130731; ROM3[6844]<=26'd9743751; ROM4[6844]<=26'd23461490;
ROM1[6845]<=26'd1956325; ROM2[6845]<=26'd11131488; ROM3[6845]<=26'd9744780; ROM4[6845]<=26'd23463318;
ROM1[6846]<=26'd1955836; ROM2[6846]<=26'd11131262; ROM3[6846]<=26'd9744524; ROM4[6846]<=26'd23463685;
ROM1[6847]<=26'd1962939; ROM2[6847]<=26'd11132445; ROM3[6847]<=26'd9741856; ROM4[6847]<=26'd23463587;
ROM1[6848]<=26'd1975428; ROM2[6848]<=26'd11135118; ROM3[6848]<=26'd9736563; ROM4[6848]<=26'd23462622;
ROM1[6849]<=26'd1977334; ROM2[6849]<=26'd11132781; ROM3[6849]<=26'd9733304; ROM4[6849]<=26'd23460016;
ROM1[6850]<=26'd1971106; ROM2[6850]<=26'd11129601; ROM3[6850]<=26'd9734772; ROM4[6850]<=26'd23459640;
ROM1[6851]<=26'd1966935; ROM2[6851]<=26'd11130694; ROM3[6851]<=26'd9739281; ROM4[6851]<=26'd23461211;
ROM1[6852]<=26'd1964142; ROM2[6852]<=26'd11133246; ROM3[6852]<=26'd9745328; ROM4[6852]<=26'd23464282;
ROM1[6853]<=26'd1960286; ROM2[6853]<=26'd11134056; ROM3[6853]<=26'd9749437; ROM4[6853]<=26'd23466368;
ROM1[6854]<=26'd1950368; ROM2[6854]<=26'd11128226; ROM3[6854]<=26'd9741287; ROM4[6854]<=26'd23457880;
ROM1[6855]<=26'd1947795; ROM2[6855]<=26'd11123444; ROM3[6855]<=26'd9733678; ROM4[6855]<=26'd23451811;
ROM1[6856]<=26'd1958344; ROM2[6856]<=26'd11121200; ROM3[6856]<=26'd9726727; ROM4[6856]<=26'd23449008;
ROM1[6857]<=26'd1969934; ROM2[6857]<=26'd11124358; ROM3[6857]<=26'd9724152; ROM4[6857]<=26'd23450535;
ROM1[6858]<=26'd1976599; ROM2[6858]<=26'd11132683; ROM3[6858]<=26'd9734201; ROM4[6858]<=26'd23459000;
ROM1[6859]<=26'd1968911; ROM2[6859]<=26'd11131290; ROM3[6859]<=26'd9736436; ROM4[6859]<=26'd23458014;
ROM1[6860]<=26'd1955579; ROM2[6860]<=26'd11124972; ROM3[6860]<=26'd9734012; ROM4[6860]<=26'd23453367;
ROM1[6861]<=26'd1948452; ROM2[6861]<=26'd11123143; ROM3[6861]<=26'd9736322; ROM4[6861]<=26'd23455059;
ROM1[6862]<=26'd1939170; ROM2[6862]<=26'd11116852; ROM3[6862]<=26'd9730824; ROM4[6862]<=26'd23449299;
ROM1[6863]<=26'd1941160; ROM2[6863]<=26'd11114820; ROM3[6863]<=26'd9727327; ROM4[6863]<=26'd23446439;
ROM1[6864]<=26'd1952999; ROM2[6864]<=26'd11115013; ROM3[6864]<=26'd9726106; ROM4[6864]<=26'd23448376;
ROM1[6865]<=26'd1966552; ROM2[6865]<=26'd11116748; ROM3[6865]<=26'd9723626; ROM4[6865]<=26'd23448979;
ROM1[6866]<=26'd1975417; ROM2[6866]<=26'd11125722; ROM3[6866]<=26'd9730979; ROM4[6866]<=26'd23457758;
ROM1[6867]<=26'd1968034; ROM2[6867]<=26'd11123912; ROM3[6867]<=26'd9731914; ROM4[6867]<=26'd23457011;
ROM1[6868]<=26'd1956139; ROM2[6868]<=26'd11117546; ROM3[6868]<=26'd9729018; ROM4[6868]<=26'd23449733;
ROM1[6869]<=26'd1948783; ROM2[6869]<=26'd11114436; ROM3[6869]<=26'd9728784; ROM4[6869]<=26'd23447839;
ROM1[6870]<=26'd1941603; ROM2[6870]<=26'd11112223; ROM3[6870]<=26'd9731887; ROM4[6870]<=26'd23448185;
ROM1[6871]<=26'd1944989; ROM2[6871]<=26'd11116187; ROM3[6871]<=26'd9735390; ROM4[6871]<=26'd23451918;
ROM1[6872]<=26'd1959927; ROM2[6872]<=26'd11125961; ROM3[6872]<=26'd9738298; ROM4[6872]<=26'd23458200;
ROM1[6873]<=26'd1980386; ROM2[6873]<=26'd11135073; ROM3[6873]<=26'd9740325; ROM4[6873]<=26'd23464509;
ROM1[6874]<=26'd1989878; ROM2[6874]<=26'd11137922; ROM3[6874]<=26'd9741357; ROM4[6874]<=26'd23466714;
ROM1[6875]<=26'd1988822; ROM2[6875]<=26'd11142110; ROM3[6875]<=26'd9747395; ROM4[6875]<=26'd23472059;
ROM1[6876]<=26'd1976432; ROM2[6876]<=26'd11137317; ROM3[6876]<=26'd9744411; ROM4[6876]<=26'd23467758;
ROM1[6877]<=26'd1966009; ROM2[6877]<=26'd11131195; ROM3[6877]<=26'd9740655; ROM4[6877]<=26'd23460359;
ROM1[6878]<=26'd1961457; ROM2[6878]<=26'd11131595; ROM3[6878]<=26'd9742905; ROM4[6878]<=26'd23460251;
ROM1[6879]<=26'd1956323; ROM2[6879]<=26'd11126143; ROM3[6879]<=26'd9741011; ROM4[6879]<=26'd23457120;
ROM1[6880]<=26'd1965197; ROM2[6880]<=26'd11128607; ROM3[6880]<=26'd9744364; ROM4[6880]<=26'd23459525;
ROM1[6881]<=26'd1981758; ROM2[6881]<=26'd11135647; ROM3[6881]<=26'd9743618; ROM4[6881]<=26'd23463861;
ROM1[6882]<=26'd1980605; ROM2[6882]<=26'd11127117; ROM3[6882]<=26'd9729233; ROM4[6882]<=26'd23454250;
ROM1[6883]<=26'd1970847; ROM2[6883]<=26'd11119632; ROM3[6883]<=26'd9720597; ROM4[6883]<=26'd23446674;
ROM1[6884]<=26'd1964798; ROM2[6884]<=26'd11120496; ROM3[6884]<=26'd9723323; ROM4[6884]<=26'd23449043;
ROM1[6885]<=26'd1954049; ROM2[6885]<=26'd11115076; ROM3[6885]<=26'd9722264; ROM4[6885]<=26'd23445895;
ROM1[6886]<=26'd1949795; ROM2[6886]<=26'd11115111; ROM3[6886]<=26'd9725503; ROM4[6886]<=26'd23447092;
ROM1[6887]<=26'd1949573; ROM2[6887]<=26'd11120735; ROM3[6887]<=26'd9731567; ROM4[6887]<=26'd23450240;
ROM1[6888]<=26'd1952329; ROM2[6888]<=26'd11121826; ROM3[6888]<=26'd9730091; ROM4[6888]<=26'd23449720;
ROM1[6889]<=26'd1966342; ROM2[6889]<=26'd11126960; ROM3[6889]<=26'd9728470; ROM4[6889]<=26'd23452195;
ROM1[6890]<=26'd1979119; ROM2[6890]<=26'd11128280; ROM3[6890]<=26'd9723945; ROM4[6890]<=26'd23452851;
ROM1[6891]<=26'd1975096; ROM2[6891]<=26'd11122994; ROM3[6891]<=26'd9720003; ROM4[6891]<=26'd23450058;
ROM1[6892]<=26'd1967107; ROM2[6892]<=26'd11121314; ROM3[6892]<=26'd9722674; ROM4[6892]<=26'd23449350;
ROM1[6893]<=26'd1961381; ROM2[6893]<=26'd11121484; ROM3[6893]<=26'd9729716; ROM4[6893]<=26'd23453226;
ROM1[6894]<=26'd1965458; ROM2[6894]<=26'd11131418; ROM3[6894]<=26'd9742100; ROM4[6894]<=26'd23463194;
ROM1[6895]<=26'd1973917; ROM2[6895]<=26'd11144194; ROM3[6895]<=26'd9755624; ROM4[6895]<=26'd23475161;
ROM1[6896]<=26'd1971492; ROM2[6896]<=26'd11140128; ROM3[6896]<=26'd9750935; ROM4[6896]<=26'd23472656;
ROM1[6897]<=26'd1967084; ROM2[6897]<=26'd11127681; ROM3[6897]<=26'd9735981; ROM4[6897]<=26'd23460711;
ROM1[6898]<=26'd1975400; ROM2[6898]<=26'd11125547; ROM3[6898]<=26'd9728389; ROM4[6898]<=26'd23457522;
ROM1[6899]<=26'd1978499; ROM2[6899]<=26'd11125296; ROM3[6899]<=26'd9723689; ROM4[6899]<=26'd23456011;
ROM1[6900]<=26'd1975769; ROM2[6900]<=26'd11127298; ROM3[6900]<=26'd9729250; ROM4[6900]<=26'd23458413;
ROM1[6901]<=26'd1974401; ROM2[6901]<=26'd11132482; ROM3[6901]<=26'd9738591; ROM4[6901]<=26'd23465123;
ROM1[6902]<=26'd1970076; ROM2[6902]<=26'd11131616; ROM3[6902]<=26'd9741250; ROM4[6902]<=26'd23467134;
ROM1[6903]<=26'd1964150; ROM2[6903]<=26'd11130764; ROM3[6903]<=26'd9745832; ROM4[6903]<=26'd23468190;
ROM1[6904]<=26'd1963781; ROM2[6904]<=26'd11131919; ROM3[6904]<=26'd9747923; ROM4[6904]<=26'd23469971;
ROM1[6905]<=26'd1966868; ROM2[6905]<=26'd11131743; ROM3[6905]<=26'd9744114; ROM4[6905]<=26'd23467762;
ROM1[6906]<=26'd1974846; ROM2[6906]<=26'd11129185; ROM3[6906]<=26'd9737256; ROM4[6906]<=26'd23463413;
ROM1[6907]<=26'd1982663; ROM2[6907]<=26'd11127259; ROM3[6907]<=26'd9733420; ROM4[6907]<=26'd23462835;
ROM1[6908]<=26'd1978175; ROM2[6908]<=26'd11125851; ROM3[6908]<=26'd9731940; ROM4[6908]<=26'd23461841;
ROM1[6909]<=26'd1971160; ROM2[6909]<=26'd11126019; ROM3[6909]<=26'd9733967; ROM4[6909]<=26'd23462454;
ROM1[6910]<=26'd1963717; ROM2[6910]<=26'd11125500; ROM3[6910]<=26'd9735398; ROM4[6910]<=26'd23459926;
ROM1[6911]<=26'd1955056; ROM2[6911]<=26'd11122743; ROM3[6911]<=26'd9734627; ROM4[6911]<=26'd23456118;
ROM1[6912]<=26'd1950258; ROM2[6912]<=26'd11122034; ROM3[6912]<=26'd9736336; ROM4[6912]<=26'd23455932;
ROM1[6913]<=26'd1953914; ROM2[6913]<=26'd11121066; ROM3[6913]<=26'd9735249; ROM4[6913]<=26'd23454901;
ROM1[6914]<=26'd1963144; ROM2[6914]<=26'd11119316; ROM3[6914]<=26'd9726618; ROM4[6914]<=26'd23451495;
ROM1[6915]<=26'd1971671; ROM2[6915]<=26'd11118685; ROM3[6915]<=26'd9718116; ROM4[6915]<=26'd23447255;
ROM1[6916]<=26'd1970069; ROM2[6916]<=26'd11117153; ROM3[6916]<=26'd9714663; ROM4[6916]<=26'd23445533;
ROM1[6917]<=26'd1962955; ROM2[6917]<=26'd11116150; ROM3[6917]<=26'd9715687; ROM4[6917]<=26'd23445208;
ROM1[6918]<=26'd1958566; ROM2[6918]<=26'd11120746; ROM3[6918]<=26'd9722388; ROM4[6918]<=26'd23449719;
ROM1[6919]<=26'd1957998; ROM2[6919]<=26'd11125090; ROM3[6919]<=26'd9729725; ROM4[6919]<=26'd23456373;
ROM1[6920]<=26'd1953331; ROM2[6920]<=26'd11123673; ROM3[6920]<=26'd9733925; ROM4[6920]<=26'd23457772;
ROM1[6921]<=26'd1953503; ROM2[6921]<=26'd11124421; ROM3[6921]<=26'd9735407; ROM4[6921]<=26'd23458791;
ROM1[6922]<=26'd1962660; ROM2[6922]<=26'd11124910; ROM3[6922]<=26'd9735137; ROM4[6922]<=26'd23461488;
ROM1[6923]<=26'd1972287; ROM2[6923]<=26'd11123360; ROM3[6923]<=26'd9725858; ROM4[6923]<=26'd23458569;
ROM1[6924]<=26'd1975524; ROM2[6924]<=26'd11123633; ROM3[6924]<=26'd9720810; ROM4[6924]<=26'd23455349;
ROM1[6925]<=26'd1967867; ROM2[6925]<=26'd11121250; ROM3[6925]<=26'd9722037; ROM4[6925]<=26'd23453322;
ROM1[6926]<=26'd1956412; ROM2[6926]<=26'd11116499; ROM3[6926]<=26'd9723418; ROM4[6926]<=26'd23450936;
ROM1[6927]<=26'd1955332; ROM2[6927]<=26'd11119132; ROM3[6927]<=26'd9732705; ROM4[6927]<=26'd23456467;
ROM1[6928]<=26'd1948620; ROM2[6928]<=26'd11119224; ROM3[6928]<=26'd9738047; ROM4[6928]<=26'd23459654;
ROM1[6929]<=26'd1943162; ROM2[6929]<=26'd11115336; ROM3[6929]<=26'd9735730; ROM4[6929]<=26'd23455757;
ROM1[6930]<=26'd1950261; ROM2[6930]<=26'd11117828; ROM3[6930]<=26'd9734793; ROM4[6930]<=26'd23456639;
ROM1[6931]<=26'd1964595; ROM2[6931]<=26'd11121671; ROM3[6931]<=26'd9732520; ROM4[6931]<=26'd23458827;
ROM1[6932]<=26'd1977224; ROM2[6932]<=26'd11125452; ROM3[6932]<=26'd9731528; ROM4[6932]<=26'd23461632;
ROM1[6933]<=26'd1976553; ROM2[6933]<=26'd11128744; ROM3[6933]<=26'd9734107; ROM4[6933]<=26'd23465573;
ROM1[6934]<=26'd1969178; ROM2[6934]<=26'd11126936; ROM3[6934]<=26'd9736865; ROM4[6934]<=26'd23463869;
ROM1[6935]<=26'd1959472; ROM2[6935]<=26'd11121915; ROM3[6935]<=26'd9735150; ROM4[6935]<=26'd23458741;
ROM1[6936]<=26'd1952146; ROM2[6936]<=26'd11120826; ROM3[6936]<=26'd9734494; ROM4[6936]<=26'd23457371;
ROM1[6937]<=26'd1946512; ROM2[6937]<=26'd11118227; ROM3[6937]<=26'd9734045; ROM4[6937]<=26'd23455416;
ROM1[6938]<=26'd1948029; ROM2[6938]<=26'd11117788; ROM3[6938]<=26'd9731066; ROM4[6938]<=26'd23454831;
ROM1[6939]<=26'd1958124; ROM2[6939]<=26'd11120328; ROM3[6939]<=26'd9726359; ROM4[6939]<=26'd23455798;
ROM1[6940]<=26'd1969752; ROM2[6940]<=26'd11120203; ROM3[6940]<=26'd9720832; ROM4[6940]<=26'd23456006;
ROM1[6941]<=26'd1974993; ROM2[6941]<=26'd11123554; ROM3[6941]<=26'd9722938; ROM4[6941]<=26'd23459435;
ROM1[6942]<=26'd1970979; ROM2[6942]<=26'd11124992; ROM3[6942]<=26'd9727521; ROM4[6942]<=26'd23461696;
ROM1[6943]<=26'd1960851; ROM2[6943]<=26'd11121835; ROM3[6943]<=26'd9729160; ROM4[6943]<=26'd23459622;
ROM1[6944]<=26'd1952041; ROM2[6944]<=26'd11118216; ROM3[6944]<=26'd9730281; ROM4[6944]<=26'd23456515;
ROM1[6945]<=26'd1945738; ROM2[6945]<=26'd11115795; ROM3[6945]<=26'd9732734; ROM4[6945]<=26'd23455781;
ROM1[6946]<=26'd1945774; ROM2[6946]<=26'd11117122; ROM3[6946]<=26'd9732888; ROM4[6946]<=26'd23457055;
ROM1[6947]<=26'd1963161; ROM2[6947]<=26'd11125739; ROM3[6947]<=26'd9738577; ROM4[6947]<=26'd23465192;
ROM1[6948]<=26'd1991211; ROM2[6948]<=26'd11141906; ROM3[6948]<=26'd9748192; ROM4[6948]<=26'd23479205;
ROM1[6949]<=26'd1991856; ROM2[6949]<=26'd11140669; ROM3[6949]<=26'd9744574; ROM4[6949]<=26'd23477404;
ROM1[6950]<=26'd1969844; ROM2[6950]<=26'd11124704; ROM3[6950]<=26'd9730100; ROM4[6950]<=26'd23461715;
ROM1[6951]<=26'd1950897; ROM2[6951]<=26'd11113307; ROM3[6951]<=26'd9720013; ROM4[6951]<=26'd23449239;
ROM1[6952]<=26'd1941101; ROM2[6952]<=26'd11108377; ROM3[6952]<=26'd9719566; ROM4[6952]<=26'd23445887;
ROM1[6953]<=26'd1935841; ROM2[6953]<=26'd11107424; ROM3[6953]<=26'd9724563; ROM4[6953]<=26'd23446842;
ROM1[6954]<=26'd1940531; ROM2[6954]<=26'd11114020; ROM3[6954]<=26'd9731869; ROM4[6954]<=26'd23453856;
ROM1[6955]<=26'd1949055; ROM2[6955]<=26'd11118112; ROM3[6955]<=26'd9735243; ROM4[6955]<=26'd23458356;
ROM1[6956]<=26'd1957033; ROM2[6956]<=26'd11115867; ROM3[6956]<=26'd9726005; ROM4[6956]<=26'd23451672;
ROM1[6957]<=26'd1966445; ROM2[6957]<=26'd11118663; ROM3[6957]<=26'd9720806; ROM4[6957]<=26'd23452244;
ROM1[6958]<=26'd1971997; ROM2[6958]<=26'd11125250; ROM3[6958]<=26'd9729860; ROM4[6958]<=26'd23459558;
ROM1[6959]<=26'd1966253; ROM2[6959]<=26'd11126482; ROM3[6959]<=26'd9735046; ROM4[6959]<=26'd23462005;
ROM1[6960]<=26'd1953448; ROM2[6960]<=26'd11119514; ROM3[6960]<=26'd9730879; ROM4[6960]<=26'd23456946;
ROM1[6961]<=26'd1945112; ROM2[6961]<=26'd11117410; ROM3[6961]<=26'd9732144; ROM4[6961]<=26'd23452982;
ROM1[6962]<=26'd1935370; ROM2[6962]<=26'd11113293; ROM3[6962]<=26'd9729468; ROM4[6962]<=26'd23448134;
ROM1[6963]<=26'd1936934; ROM2[6963]<=26'd11111308; ROM3[6963]<=26'd9725297; ROM4[6963]<=26'd23445316;
ROM1[6964]<=26'd1951186; ROM2[6964]<=26'd11115821; ROM3[6964]<=26'd9724272; ROM4[6964]<=26'd23448081;
ROM1[6965]<=26'd1965111; ROM2[6965]<=26'd11118445; ROM3[6965]<=26'd9718749; ROM4[6965]<=26'd23448218;
ROM1[6966]<=26'd1965602; ROM2[6966]<=26'd11118530; ROM3[6966]<=26'd9716562; ROM4[6966]<=26'd23446056;
ROM1[6967]<=26'd1957100; ROM2[6967]<=26'd11116075; ROM3[6967]<=26'd9716858; ROM4[6967]<=26'd23444768;
ROM1[6968]<=26'd1949368; ROM2[6968]<=26'd11114173; ROM3[6968]<=26'd9721417; ROM4[6968]<=26'd23445669;
ROM1[6969]<=26'd1942044; ROM2[6969]<=26'd11113012; ROM3[6969]<=26'd9725148; ROM4[6969]<=26'd23446938;
ROM1[6970]<=26'd1936385; ROM2[6970]<=26'd11111644; ROM3[6970]<=26'd9728449; ROM4[6970]<=26'd23447414;
ROM1[6971]<=26'd1937530; ROM2[6971]<=26'd11111421; ROM3[6971]<=26'd9730796; ROM4[6971]<=26'd23447191;
ROM1[6972]<=26'd1946094; ROM2[6972]<=26'd11113001; ROM3[6972]<=26'd9729051; ROM4[6972]<=26'd23445573;
ROM1[6973]<=26'd1960239; ROM2[6973]<=26'd11114997; ROM3[6973]<=26'd9723084; ROM4[6973]<=26'd23445615;
ROM1[6974]<=26'd1965198; ROM2[6974]<=26'd11115443; ROM3[6974]<=26'd9720259; ROM4[6974]<=26'd23446373;
ROM1[6975]<=26'd1960677; ROM2[6975]<=26'd11116656; ROM3[6975]<=26'd9725535; ROM4[6975]<=26'd23448782;
ROM1[6976]<=26'd1953535; ROM2[6976]<=26'd11114335; ROM3[6976]<=26'd9729067; ROM4[6976]<=26'd23450330;
ROM1[6977]<=26'd1948720; ROM2[6977]<=26'd11111592; ROM3[6977]<=26'd9732410; ROM4[6977]<=26'd23450053;
ROM1[6978]<=26'd1944783; ROM2[6978]<=26'd11113468; ROM3[6978]<=26'd9738112; ROM4[6978]<=26'd23452109;
ROM1[6979]<=26'd1938021; ROM2[6979]<=26'd11109482; ROM3[6979]<=26'd9734409; ROM4[6979]<=26'd23448205;
ROM1[6980]<=26'd1945085; ROM2[6980]<=26'd11111270; ROM3[6980]<=26'd9733006; ROM4[6980]<=26'd23449226;
ROM1[6981]<=26'd1960958; ROM2[6981]<=26'd11117955; ROM3[6981]<=26'd9733160; ROM4[6981]<=26'd23455794;
ROM1[6982]<=26'd1968366; ROM2[6982]<=26'd11119236; ROM3[6982]<=26'd9729851; ROM4[6982]<=26'd23457205;
ROM1[6983]<=26'd1963124; ROM2[6983]<=26'd11113923; ROM3[6983]<=26'd9728333; ROM4[6983]<=26'd23454874;
ROM1[6984]<=26'd1954417; ROM2[6984]<=26'd11111635; ROM3[6984]<=26'd9729282; ROM4[6984]<=26'd23452525;
ROM1[6985]<=26'd1950459; ROM2[6985]<=26'd11113089; ROM3[6985]<=26'd9731607; ROM4[6985]<=26'd23452760;
ROM1[6986]<=26'd1943865; ROM2[6986]<=26'd11111622; ROM3[6986]<=26'd9731956; ROM4[6986]<=26'd23451700;
ROM1[6987]<=26'd1939640; ROM2[6987]<=26'd11113331; ROM3[6987]<=26'd9733263; ROM4[6987]<=26'd23451387;
ROM1[6988]<=26'd1941370; ROM2[6988]<=26'd11113607; ROM3[6988]<=26'd9730372; ROM4[6988]<=26'd23450446;
ROM1[6989]<=26'd1946945; ROM2[6989]<=26'd11111091; ROM3[6989]<=26'd9723077; ROM4[6989]<=26'd23446363;
ROM1[6990]<=26'd1959658; ROM2[6990]<=26'd11113461; ROM3[6990]<=26'd9720959; ROM4[6990]<=26'd23446947;
ROM1[6991]<=26'd1965995; ROM2[6991]<=26'd11119882; ROM3[6991]<=26'd9725009; ROM4[6991]<=26'd23452507;
ROM1[6992]<=26'd1962462; ROM2[6992]<=26'd11122068; ROM3[6992]<=26'd9730225; ROM4[6992]<=26'd23455349;
ROM1[6993]<=26'd1955249; ROM2[6993]<=26'd11120136; ROM3[6993]<=26'd9735775; ROM4[6993]<=26'd23454376;
ROM1[6994]<=26'd1952305; ROM2[6994]<=26'd11121495; ROM3[6994]<=26'd9739488; ROM4[6994]<=26'd23457720;
ROM1[6995]<=26'd1952193; ROM2[6995]<=26'd11125540; ROM3[6995]<=26'd9746237; ROM4[6995]<=26'd23463168;
ROM1[6996]<=26'd1949382; ROM2[6996]<=26'd11122088; ROM3[6996]<=26'd9742569; ROM4[6996]<=26'd23460181;
ROM1[6997]<=26'd1952383; ROM2[6997]<=26'd11118543; ROM3[6997]<=26'd9732731; ROM4[6997]<=26'd23455869;
ROM1[6998]<=26'd1968092; ROM2[6998]<=26'd11121830; ROM3[6998]<=26'd9730399; ROM4[6998]<=26'd23456488;
ROM1[6999]<=26'd1970585; ROM2[6999]<=26'd11119805; ROM3[6999]<=26'd9726944; ROM4[6999]<=26'd23454634;
ROM1[7000]<=26'd1960374; ROM2[7000]<=26'd11116224; ROM3[7000]<=26'd9725485; ROM4[7000]<=26'd23451368;
ROM1[7001]<=26'd1961700; ROM2[7001]<=26'd11125051; ROM3[7001]<=26'd9736842; ROM4[7001]<=26'd23459679;
ROM1[7002]<=26'd1954609; ROM2[7002]<=26'd11121341; ROM3[7002]<=26'd9736484; ROM4[7002]<=26'd23456429;
ROM1[7003]<=26'd1939203; ROM2[7003]<=26'd11109596; ROM3[7003]<=26'd9728034; ROM4[7003]<=26'd23445521;
ROM1[7004]<=26'd1937359; ROM2[7004]<=26'd11109777; ROM3[7004]<=26'd9729026; ROM4[7004]<=26'd23446424;
ROM1[7005]<=26'd1946915; ROM2[7005]<=26'd11114136; ROM3[7005]<=26'd9731397; ROM4[7005]<=26'd23449570;
ROM1[7006]<=26'd1967979; ROM2[7006]<=26'd11123411; ROM3[7006]<=26'd9733272; ROM4[7006]<=26'd23456503;
ROM1[7007]<=26'd1980858; ROM2[7007]<=26'd11128884; ROM3[7007]<=26'd9732284; ROM4[7007]<=26'd23460387;
ROM1[7008]<=26'd1972966; ROM2[7008]<=26'd11123475; ROM3[7008]<=26'd9729241; ROM4[7008]<=26'd23454981;
ROM1[7009]<=26'd1957626; ROM2[7009]<=26'd11114123; ROM3[7009]<=26'd9724774; ROM4[7009]<=26'd23447282;
ROM1[7010]<=26'd1946581; ROM2[7010]<=26'd11108826; ROM3[7010]<=26'd9724686; ROM4[7010]<=26'd23444757;
ROM1[7011]<=26'd1944240; ROM2[7011]<=26'd11110641; ROM3[7011]<=26'd9731358; ROM4[7011]<=26'd23446848;
ROM1[7012]<=26'd1946538; ROM2[7012]<=26'd11118073; ROM3[7012]<=26'd9737704; ROM4[7012]<=26'd23452808;
ROM1[7013]<=26'd1951436; ROM2[7013]<=26'd11121209; ROM3[7013]<=26'd9739003; ROM4[7013]<=26'd23456353;
ROM1[7014]<=26'd1960710; ROM2[7014]<=26'd11120447; ROM3[7014]<=26'd9734078; ROM4[7014]<=26'd23453603;
ROM1[7015]<=26'd1972445; ROM2[7015]<=26'd11123556; ROM3[7015]<=26'd9731245; ROM4[7015]<=26'd23454253;
ROM1[7016]<=26'd1974563; ROM2[7016]<=26'd11124448; ROM3[7016]<=26'd9732747; ROM4[7016]<=26'd23456512;
ROM1[7017]<=26'd1967824; ROM2[7017]<=26'd11121614; ROM3[7017]<=26'd9734569; ROM4[7017]<=26'd23456301;
ROM1[7018]<=26'd1958373; ROM2[7018]<=26'd11118727; ROM3[7018]<=26'd9734942; ROM4[7018]<=26'd23455016;
ROM1[7019]<=26'd1951491; ROM2[7019]<=26'd11117199; ROM3[7019]<=26'd9735025; ROM4[7019]<=26'd23455429;
ROM1[7020]<=26'd1947358; ROM2[7020]<=26'd11118671; ROM3[7020]<=26'd9739704; ROM4[7020]<=26'd23457496;
ROM1[7021]<=26'd1948442; ROM2[7021]<=26'd11119185; ROM3[7021]<=26'd9738453; ROM4[7021]<=26'd23457392;
ROM1[7022]<=26'd1958445; ROM2[7022]<=26'd11121586; ROM3[7022]<=26'd9734565; ROM4[7022]<=26'd23457161;
ROM1[7023]<=26'd1970243; ROM2[7023]<=26'd11121381; ROM3[7023]<=26'd9726069; ROM4[7023]<=26'd23454733;
ROM1[7024]<=26'd1972087; ROM2[7024]<=26'd11117836; ROM3[7024]<=26'd9721133; ROM4[7024]<=26'd23451968;
ROM1[7025]<=26'd1966932; ROM2[7025]<=26'd11118213; ROM3[7025]<=26'd9721935; ROM4[7025]<=26'd23450554;
ROM1[7026]<=26'd1962008; ROM2[7026]<=26'd11120998; ROM3[7026]<=26'd9727150; ROM4[7026]<=26'd23453031;
ROM1[7027]<=26'd1962041; ROM2[7027]<=26'd11124979; ROM3[7027]<=26'd9736600; ROM4[7027]<=26'd23459008;
ROM1[7028]<=26'd1958336; ROM2[7028]<=26'd11126238; ROM3[7028]<=26'd9740666; ROM4[7028]<=26'd23460481;
ROM1[7029]<=26'd1952864; ROM2[7029]<=26'd11124182; ROM3[7029]<=26'd9740046; ROM4[7029]<=26'd23459685;
ROM1[7030]<=26'd1957842; ROM2[7030]<=26'd11125518; ROM3[7030]<=26'd9739357; ROM4[7030]<=26'd23459277;
ROM1[7031]<=26'd1972638; ROM2[7031]<=26'd11129169; ROM3[7031]<=26'd9736284; ROM4[7031]<=26'd23459461;
ROM1[7032]<=26'd1981611; ROM2[7032]<=26'd11129120; ROM3[7032]<=26'd9733557; ROM4[7032]<=26'd23459085;
ROM1[7033]<=26'd1980602; ROM2[7033]<=26'd11131345; ROM3[7033]<=26'd9739405; ROM4[7033]<=26'd23462452;
ROM1[7034]<=26'd1970925; ROM2[7034]<=26'd11127182; ROM3[7034]<=26'd9741752; ROM4[7034]<=26'd23461504;
ROM1[7035]<=26'd1959502; ROM2[7035]<=26'd11120175; ROM3[7035]<=26'd9740052; ROM4[7035]<=26'd23455447;
ROM1[7036]<=26'd1953189; ROM2[7036]<=26'd11120161; ROM3[7036]<=26'd9740957; ROM4[7036]<=26'd23455675;
ROM1[7037]<=26'd1953543; ROM2[7037]<=26'd11123724; ROM3[7037]<=26'd9746816; ROM4[7037]<=26'd23460176;
ROM1[7038]<=26'd1962547; ROM2[7038]<=26'd11130737; ROM3[7038]<=26'd9751793; ROM4[7038]<=26'd23466058;
ROM1[7039]<=26'd1973715; ROM2[7039]<=26'd11134223; ROM3[7039]<=26'd9747424; ROM4[7039]<=26'd23466808;
ROM1[7040]<=26'd1984911; ROM2[7040]<=26'd11133695; ROM3[7040]<=26'd9741445; ROM4[7040]<=26'd23465219;
ROM1[7041]<=26'd1975006; ROM2[7041]<=26'd11121100; ROM3[7041]<=26'd9729178; ROM4[7041]<=26'd23455650;
ROM1[7042]<=26'd1964880; ROM2[7042]<=26'd11117380; ROM3[7042]<=26'd9727506; ROM4[7042]<=26'd23454219;
ROM1[7043]<=26'd1961234; ROM2[7043]<=26'd11121567; ROM3[7043]<=26'd9734739; ROM4[7043]<=26'd23458902;
ROM1[7044]<=26'd1958290; ROM2[7044]<=26'd11124292; ROM3[7044]<=26'd9738936; ROM4[7044]<=26'd23461999;
ROM1[7045]<=26'd1960663; ROM2[7045]<=26'd11131914; ROM3[7045]<=26'd9746665; ROM4[7045]<=26'd23467646;
ROM1[7046]<=26'd1958847; ROM2[7046]<=26'd11128987; ROM3[7046]<=26'd9744907; ROM4[7046]<=26'd23463666;
ROM1[7047]<=26'd1960840; ROM2[7047]<=26'd11122935; ROM3[7047]<=26'd9737017; ROM4[7047]<=26'd23458586;
ROM1[7048]<=26'd1971429; ROM2[7048]<=26'd11122315; ROM3[7048]<=26'd9731324; ROM4[7048]<=26'd23457179;
ROM1[7049]<=26'd1976396; ROM2[7049]<=26'd11124168; ROM3[7049]<=26'd9728605; ROM4[7049]<=26'd23456610;
ROM1[7050]<=26'd1973135; ROM2[7050]<=26'd11125590; ROM3[7050]<=26'd9731337; ROM4[7050]<=26'd23458299;
ROM1[7051]<=26'd1968053; ROM2[7051]<=26'd11125914; ROM3[7051]<=26'd9736206; ROM4[7051]<=26'd23460045;
ROM1[7052]<=26'd1963773; ROM2[7052]<=26'd11125717; ROM3[7052]<=26'd9739155; ROM4[7052]<=26'd23461152;
ROM1[7053]<=26'd1956659; ROM2[7053]<=26'd11123683; ROM3[7053]<=26'd9742569; ROM4[7053]<=26'd23461213;
ROM1[7054]<=26'd1953219; ROM2[7054]<=26'd11121806; ROM3[7054]<=26'd9741724; ROM4[7054]<=26'd23460554;
ROM1[7055]<=26'd1959404; ROM2[7055]<=26'd11122225; ROM3[7055]<=26'd9738602; ROM4[7055]<=26'd23459557;
ROM1[7056]<=26'd1973927; ROM2[7056]<=26'd11124584; ROM3[7056]<=26'd9733878; ROM4[7056]<=26'd23458819;
ROM1[7057]<=26'd1983578; ROM2[7057]<=26'd11126763; ROM3[7057]<=26'd9732612; ROM4[7057]<=26'd23459350;
ROM1[7058]<=26'd1981404; ROM2[7058]<=26'd11128941; ROM3[7058]<=26'd9737104; ROM4[7058]<=26'd23461737;
ROM1[7059]<=26'd1972509; ROM2[7059]<=26'd11127331; ROM3[7059]<=26'd9740377; ROM4[7059]<=26'd23461128;
ROM1[7060]<=26'd1966018; ROM2[7060]<=26'd11125415; ROM3[7060]<=26'd9745983; ROM4[7060]<=26'd23461814;
ROM1[7061]<=26'd1963328; ROM2[7061]<=26'd11125449; ROM3[7061]<=26'd9752609; ROM4[7061]<=26'd23465696;
ROM1[7062]<=26'd1951972; ROM2[7062]<=26'd11118149; ROM3[7062]<=26'd9749089; ROM4[7062]<=26'd23460488;
ROM1[7063]<=26'd1951884; ROM2[7063]<=26'd11117555; ROM3[7063]<=26'd9747308; ROM4[7063]<=26'd23459278;
ROM1[7064]<=26'd1965000; ROM2[7064]<=26'd11123450; ROM3[7064]<=26'd9740974; ROM4[7064]<=26'd23458035;
ROM1[7065]<=26'd1978785; ROM2[7065]<=26'd11126493; ROM3[7065]<=26'd9732448; ROM4[7065]<=26'd23455616;
ROM1[7066]<=26'd1983948; ROM2[7066]<=26'd11129645; ROM3[7066]<=26'd9735220; ROM4[7066]<=26'd23458447;
ROM1[7067]<=26'd1977645; ROM2[7067]<=26'd11129345; ROM3[7067]<=26'd9737315; ROM4[7067]<=26'd23460735;
ROM1[7068]<=26'd1969367; ROM2[7068]<=26'd11128254; ROM3[7068]<=26'd9739913; ROM4[7068]<=26'd23461052;
ROM1[7069]<=26'd1961968; ROM2[7069]<=26'd11127352; ROM3[7069]<=26'd9740150; ROM4[7069]<=26'd23458957;
ROM1[7070]<=26'd1955813; ROM2[7070]<=26'd11124355; ROM3[7070]<=26'd9739080; ROM4[7070]<=26'd23456375;
ROM1[7071]<=26'd1958422; ROM2[7071]<=26'd11123701; ROM3[7071]<=26'd9739793; ROM4[7071]<=26'd23455274;
ROM1[7072]<=26'd1966486; ROM2[7072]<=26'd11124799; ROM3[7072]<=26'd9738686; ROM4[7072]<=26'd23456408;
ROM1[7073]<=26'd1978344; ROM2[7073]<=26'd11125857; ROM3[7073]<=26'd9733988; ROM4[7073]<=26'd23458469;
ROM1[7074]<=26'd1989723; ROM2[7074]<=26'd11134026; ROM3[7074]<=26'd9740381; ROM4[7074]<=26'd23467968;
ROM1[7075]<=26'd1988474; ROM2[7075]<=26'd11137662; ROM3[7075]<=26'd9745611; ROM4[7075]<=26'd23472302;
ROM1[7076]<=26'd1970965; ROM2[7076]<=26'd11127105; ROM3[7076]<=26'd9740414; ROM4[7076]<=26'd23463956;
ROM1[7077]<=26'd1958529; ROM2[7077]<=26'd11120823; ROM3[7077]<=26'd9738514; ROM4[7077]<=26'd23458843;
ROM1[7078]<=26'd1953094; ROM2[7078]<=26'd11120715; ROM3[7078]<=26'd9740209; ROM4[7078]<=26'd23457963;
ROM1[7079]<=26'd1952493; ROM2[7079]<=26'd11120758; ROM3[7079]<=26'd9744919; ROM4[7079]<=26'd23460708;
ROM1[7080]<=26'd1964095; ROM2[7080]<=26'd11126987; ROM3[7080]<=26'd9751001; ROM4[7080]<=26'd23467579;
ROM1[7081]<=26'd1975775; ROM2[7081]<=26'd11127248; ROM3[7081]<=26'd9746000; ROM4[7081]<=26'd23465890;
ROM1[7082]<=26'd1978606; ROM2[7082]<=26'd11120942; ROM3[7082]<=26'd9736125; ROM4[7082]<=26'd23459170;
ROM1[7083]<=26'd1970942; ROM2[7083]<=26'd11116614; ROM3[7083]<=26'd9731043; ROM4[7083]<=26'd23454858;
ROM1[7084]<=26'd1961569; ROM2[7084]<=26'd11115547; ROM3[7084]<=26'd9731595; ROM4[7084]<=26'd23453118;
ROM1[7085]<=26'd1958530; ROM2[7085]<=26'd11116554; ROM3[7085]<=26'd9737640; ROM4[7085]<=26'd23454248;
ROM1[7086]<=26'd1956410; ROM2[7086]<=26'd11118957; ROM3[7086]<=26'd9742844; ROM4[7086]<=26'd23457483;
ROM1[7087]<=26'd1960647; ROM2[7087]<=26'd11128327; ROM3[7087]<=26'd9750310; ROM4[7087]<=26'd23464779;
ROM1[7088]<=26'd1969277; ROM2[7088]<=26'd11132552; ROM3[7088]<=26'd9753373; ROM4[7088]<=26'd23468730;
ROM1[7089]<=26'd1972206; ROM2[7089]<=26'd11125548; ROM3[7089]<=26'd9740581; ROM4[7089]<=26'd23460336;
ROM1[7090]<=26'd1974581; ROM2[7090]<=26'd11118431; ROM3[7090]<=26'd9727039; ROM4[7090]<=26'd23449803;
ROM1[7091]<=26'd1971023; ROM2[7091]<=26'd11115647; ROM3[7091]<=26'd9723796; ROM4[7091]<=26'd23446616;
ROM1[7092]<=26'd1964067; ROM2[7092]<=26'd11115502; ROM3[7092]<=26'd9725542; ROM4[7092]<=26'd23447915;
ROM1[7093]<=26'd1957780; ROM2[7093]<=26'd11116542; ROM3[7093]<=26'd9729353; ROM4[7093]<=26'd23450691;
ROM1[7094]<=26'd1950650; ROM2[7094]<=26'd11114533; ROM3[7094]<=26'd9730305; ROM4[7094]<=26'd23451225;
ROM1[7095]<=26'd1940557; ROM2[7095]<=26'd11107987; ROM3[7095]<=26'd9727661; ROM4[7095]<=26'd23447087;
ROM1[7096]<=26'd1938750; ROM2[7096]<=26'd11104916; ROM3[7096]<=26'd9724767; ROM4[7096]<=26'd23444933;
ROM1[7097]<=26'd1950337; ROM2[7097]<=26'd11109085; ROM3[7097]<=26'd9724856; ROM4[7097]<=26'd23448898;
ROM1[7098]<=26'd1967040; ROM2[7098]<=26'd11114581; ROM3[7098]<=26'd9723955; ROM4[7098]<=26'd23452864;
ROM1[7099]<=26'd1973130; ROM2[7099]<=26'd11117181; ROM3[7099]<=26'd9724763; ROM4[7099]<=26'd23454811;
ROM1[7100]<=26'd1967084; ROM2[7100]<=26'd11116220; ROM3[7100]<=26'd9726200; ROM4[7100]<=26'd23453186;
ROM1[7101]<=26'd1963418; ROM2[7101]<=26'd11118424; ROM3[7101]<=26'd9731791; ROM4[7101]<=26'd23454673;
ROM1[7102]<=26'd1961537; ROM2[7102]<=26'd11123323; ROM3[7102]<=26'd9738159; ROM4[7102]<=26'd23459856;
ROM1[7103]<=26'd1957146; ROM2[7103]<=26'd11123672; ROM3[7103]<=26'd9740888; ROM4[7103]<=26'd23459931;
ROM1[7104]<=26'd1957324; ROM2[7104]<=26'd11124862; ROM3[7104]<=26'd9743956; ROM4[7104]<=26'd23462274;
ROM1[7105]<=26'd1960195; ROM2[7105]<=26'd11123618; ROM3[7105]<=26'd9742399; ROM4[7105]<=26'd23461296;
ROM1[7106]<=26'd1969932; ROM2[7106]<=26'd11121171; ROM3[7106]<=26'd9736941; ROM4[7106]<=26'd23457112;
ROM1[7107]<=26'd1974844; ROM2[7107]<=26'd11119911; ROM3[7107]<=26'd9732048; ROM4[7107]<=26'd23455781;
ROM1[7108]<=26'd1970516; ROM2[7108]<=26'd11118918; ROM3[7108]<=26'd9732818; ROM4[7108]<=26'd23456376;
ROM1[7109]<=26'd1969569; ROM2[7109]<=26'd11123194; ROM3[7109]<=26'd9740730; ROM4[7109]<=26'd23461365;
ROM1[7110]<=26'd1965348; ROM2[7110]<=26'd11123624; ROM3[7110]<=26'd9743697; ROM4[7110]<=26'd23462499;
ROM1[7111]<=26'd1959294; ROM2[7111]<=26'd11120791; ROM3[7111]<=26'd9745352; ROM4[7111]<=26'd23461618;
ROM1[7112]<=26'd1956096; ROM2[7112]<=26'd11122165; ROM3[7112]<=26'd9746928; ROM4[7112]<=26'd23463241;
ROM1[7113]<=26'd1958271; ROM2[7113]<=26'd11124029; ROM3[7113]<=26'd9746235; ROM4[7113]<=26'd23465064;
ROM1[7114]<=26'd1972815; ROM2[7114]<=26'd11130221; ROM3[7114]<=26'd9746180; ROM4[7114]<=26'd23468072;
ROM1[7115]<=26'd1986045; ROM2[7115]<=26'd11133920; ROM3[7115]<=26'd9744265; ROM4[7115]<=26'd23470951;
ROM1[7116]<=26'd1982507; ROM2[7116]<=26'd11128796; ROM3[7116]<=26'd9742645; ROM4[7116]<=26'd23467680;
ROM1[7117]<=26'd1973687; ROM2[7117]<=26'd11124024; ROM3[7117]<=26'd9740553; ROM4[7117]<=26'd23463709;
ROM1[7118]<=26'd1966602; ROM2[7118]<=26'd11124494; ROM3[7118]<=26'd9744190; ROM4[7118]<=26'd23465400;
ROM1[7119]<=26'd1963461; ROM2[7119]<=26'd11127491; ROM3[7119]<=26'd9749465; ROM4[7119]<=26'd23468098;
ROM1[7120]<=26'd1956744; ROM2[7120]<=26'd11124712; ROM3[7120]<=26'd9747289; ROM4[7120]<=26'd23464307;
ROM1[7121]<=26'd1955324; ROM2[7121]<=26'd11122314; ROM3[7121]<=26'd9745588; ROM4[7121]<=26'd23460884;
ROM1[7122]<=26'd1963082; ROM2[7122]<=26'd11120897; ROM3[7122]<=26'd9741932; ROM4[7122]<=26'd23460030;
ROM1[7123]<=26'd1974638; ROM2[7123]<=26'd11120167; ROM3[7123]<=26'd9736047; ROM4[7123]<=26'd23458333;
ROM1[7124]<=26'd1980579; ROM2[7124]<=26'd11122160; ROM3[7124]<=26'd9737096; ROM4[7124]<=26'd23460501;
ROM1[7125]<=26'd1974521; ROM2[7125]<=26'd11120742; ROM3[7125]<=26'd9738137; ROM4[7125]<=26'd23461188;
ROM1[7126]<=26'd1966045; ROM2[7126]<=26'd11117406; ROM3[7126]<=26'd9738807; ROM4[7126]<=26'd23459971;
ROM1[7127]<=26'd1969777; ROM2[7127]<=26'd11124432; ROM3[7127]<=26'd9747418; ROM4[7127]<=26'd23468165;
ROM1[7128]<=26'd1969374; ROM2[7128]<=26'd11129789; ROM3[7128]<=26'd9754626; ROM4[7128]<=26'd23474437;
ROM1[7129]<=26'd1967464; ROM2[7129]<=26'd11130584; ROM3[7129]<=26'd9756388; ROM4[7129]<=26'd23476075;
ROM1[7130]<=26'd1967767; ROM2[7130]<=26'd11127390; ROM3[7130]<=26'd9750653; ROM4[7130]<=26'd23471688;
ROM1[7131]<=26'd1972191; ROM2[7131]<=26'd11120302; ROM3[7131]<=26'd9736109; ROM4[7131]<=26'd23461685;
ROM1[7132]<=26'd1984294; ROM2[7132]<=26'd11123357; ROM3[7132]<=26'd9732616; ROM4[7132]<=26'd23462101;
ROM1[7133]<=26'd1983548; ROM2[7133]<=26'd11126941; ROM3[7133]<=26'd9734463; ROM4[7133]<=26'd23463612;
ROM1[7134]<=26'd1975436; ROM2[7134]<=26'd11126515; ROM3[7134]<=26'd9736153; ROM4[7134]<=26'd23463517;
ROM1[7135]<=26'd1969544; ROM2[7135]<=26'd11126079; ROM3[7135]<=26'd9741069; ROM4[7135]<=26'd23465440;
ROM1[7136]<=26'd1961362; ROM2[7136]<=26'd11122477; ROM3[7136]<=26'd9739701; ROM4[7136]<=26'd23462390;
ROM1[7137]<=26'd1956537; ROM2[7137]<=26'd11121138; ROM3[7137]<=26'd9739913; ROM4[7137]<=26'd23459371;
ROM1[7138]<=26'd1961436; ROM2[7138]<=26'd11124203; ROM3[7138]<=26'd9739121; ROM4[7138]<=26'd23460296;
ROM1[7139]<=26'd1973722; ROM2[7139]<=26'd11129241; ROM3[7139]<=26'd9734709; ROM4[7139]<=26'd23461365;
ROM1[7140]<=26'd1981771; ROM2[7140]<=26'd11128177; ROM3[7140]<=26'd9730296; ROM4[7140]<=26'd23459573;
ROM1[7141]<=26'd1974253; ROM2[7141]<=26'd11119132; ROM3[7141]<=26'd9723526; ROM4[7141]<=26'd23453313;
ROM1[7142]<=26'd1966641; ROM2[7142]<=26'd11116990; ROM3[7142]<=26'd9725447; ROM4[7142]<=26'd23452120;
ROM1[7143]<=26'd1955825; ROM2[7143]<=26'd11112215; ROM3[7143]<=26'd9727346; ROM4[7143]<=26'd23449558;
ROM1[7144]<=26'd1948222; ROM2[7144]<=26'd11109310; ROM3[7144]<=26'd9728148; ROM4[7144]<=26'd23448805;
ROM1[7145]<=26'd1948943; ROM2[7145]<=26'd11113967; ROM3[7145]<=26'd9735270; ROM4[7145]<=26'd23454208;
ROM1[7146]<=26'd1951292; ROM2[7146]<=26'd11114326; ROM3[7146]<=26'd9736278; ROM4[7146]<=26'd23453898;
ROM1[7147]<=26'd1958326; ROM2[7147]<=26'd11112071; ROM3[7147]<=26'd9730351; ROM4[7147]<=26'd23450617;
ROM1[7148]<=26'd1968096; ROM2[7148]<=26'd11110774; ROM3[7148]<=26'd9723127; ROM4[7148]<=26'd23445665;
ROM1[7149]<=26'd1973589; ROM2[7149]<=26'd11113865; ROM3[7149]<=26'd9724547; ROM4[7149]<=26'd23449734;
ROM1[7150]<=26'd1969797; ROM2[7150]<=26'd11114752; ROM3[7150]<=26'd9729471; ROM4[7150]<=26'd23453466;
ROM1[7151]<=26'd1964566; ROM2[7151]<=26'd11117027; ROM3[7151]<=26'd9736968; ROM4[7151]<=26'd23455328;
ROM1[7152]<=26'd1966281; ROM2[7152]<=26'd11124368; ROM3[7152]<=26'd9746135; ROM4[7152]<=26'd23463171;
ROM1[7153]<=26'd1965194; ROM2[7153]<=26'd11126853; ROM3[7153]<=26'd9750141; ROM4[7153]<=26'd23464448;
ROM1[7154]<=26'd1957989; ROM2[7154]<=26'd11118825; ROM3[7154]<=26'd9742156; ROM4[7154]<=26'd23456525;
ROM1[7155]<=26'd1958368; ROM2[7155]<=26'd11114835; ROM3[7155]<=26'd9734095; ROM4[7155]<=26'd23450893;
ROM1[7156]<=26'd1970724; ROM2[7156]<=26'd11119591; ROM3[7156]<=26'd9730885; ROM4[7156]<=26'd23451757;
ROM1[7157]<=26'd1974040; ROM2[7157]<=26'd11118032; ROM3[7157]<=26'd9723657; ROM4[7157]<=26'd23449211;
ROM1[7158]<=26'd1970325; ROM2[7158]<=26'd11117756; ROM3[7158]<=26'd9726543; ROM4[7158]<=26'd23449843;
ROM1[7159]<=26'd1965486; ROM2[7159]<=26'd11119672; ROM3[7159]<=26'd9730777; ROM4[7159]<=26'd23451326;
ROM1[7160]<=26'd1958530; ROM2[7160]<=26'd11115829; ROM3[7160]<=26'd9730137; ROM4[7160]<=26'd23448406;
ROM1[7161]<=26'd1954812; ROM2[7161]<=26'd11116025; ROM3[7161]<=26'd9736528; ROM4[7161]<=26'd23450626;
ROM1[7162]<=26'd1952434; ROM2[7162]<=26'd11120007; ROM3[7162]<=26'd9739332; ROM4[7162]<=26'd23454258;
ROM1[7163]<=26'd1955843; ROM2[7163]<=26'd11120422; ROM3[7163]<=26'd9737871; ROM4[7163]<=26'd23454849;
ROM1[7164]<=26'd1965435; ROM2[7164]<=26'd11120402; ROM3[7164]<=26'd9734101; ROM4[7164]<=26'd23454562;
ROM1[7165]<=26'd1976444; ROM2[7165]<=26'd11120221; ROM3[7165]<=26'd9729125; ROM4[7165]<=26'd23455008;
ROM1[7166]<=26'd1979844; ROM2[7166]<=26'd11123268; ROM3[7166]<=26'd9734034; ROM4[7166]<=26'd23458234;
ROM1[7167]<=26'd1975809; ROM2[7167]<=26'd11126445; ROM3[7167]<=26'd9740583; ROM4[7167]<=26'd23462304;
ROM1[7168]<=26'd1967685; ROM2[7168]<=26'd11126466; ROM3[7168]<=26'd9744604; ROM4[7168]<=26'd23464500;
ROM1[7169]<=26'd1960674; ROM2[7169]<=26'd11123836; ROM3[7169]<=26'd9747056; ROM4[7169]<=26'd23463405;
ROM1[7170]<=26'd1952340; ROM2[7170]<=26'd11120080; ROM3[7170]<=26'd9745775; ROM4[7170]<=26'd23460372;
ROM1[7171]<=26'd1949280; ROM2[7171]<=26'd11115754; ROM3[7171]<=26'd9741810; ROM4[7171]<=26'd23456725;
ROM1[7172]<=26'd1957238; ROM2[7172]<=26'd11112787; ROM3[7172]<=26'd9737857; ROM4[7172]<=26'd23454413;
ROM1[7173]<=26'd1967402; ROM2[7173]<=26'd11113860; ROM3[7173]<=26'd9731590; ROM4[7173]<=26'd23453872;
ROM1[7174]<=26'd1967643; ROM2[7174]<=26'd11113569; ROM3[7174]<=26'd9727829; ROM4[7174]<=26'd23450708;
ROM1[7175]<=26'd1961911; ROM2[7175]<=26'd11112910; ROM3[7175]<=26'd9730377; ROM4[7175]<=26'd23449971;
ROM1[7176]<=26'd1956928; ROM2[7176]<=26'd11114386; ROM3[7176]<=26'd9734114; ROM4[7176]<=26'd23451085;
ROM1[7177]<=26'd1952319; ROM2[7177]<=26'd11114969; ROM3[7177]<=26'd9736537; ROM4[7177]<=26'd23451374;
ROM1[7178]<=26'd1946371; ROM2[7178]<=26'd11114748; ROM3[7178]<=26'd9741137; ROM4[7178]<=26'd23453829;
ROM1[7179]<=26'd1947290; ROM2[7179]<=26'd11118281; ROM3[7179]<=26'd9744852; ROM4[7179]<=26'd23456998;
ROM1[7180]<=26'd1952838; ROM2[7180]<=26'd11120056; ROM3[7180]<=26'd9743255; ROM4[7180]<=26'd23456355;
ROM1[7181]<=26'd1965973; ROM2[7181]<=26'd11121924; ROM3[7181]<=26'd9738353; ROM4[7181]<=26'd23455705;
ROM1[7182]<=26'd1976843; ROM2[7182]<=26'd11122504; ROM3[7182]<=26'd9735097; ROM4[7182]<=26'd23454329;
ROM1[7183]<=26'd1970307; ROM2[7183]<=26'd11118332; ROM3[7183]<=26'd9733625; ROM4[7183]<=26'd23451453;
ROM1[7184]<=26'd1959775; ROM2[7184]<=26'd11115660; ROM3[7184]<=26'd9735305; ROM4[7184]<=26'd23450874;
ROM1[7185]<=26'd1954151; ROM2[7185]<=26'd11115513; ROM3[7185]<=26'd9739793; ROM4[7185]<=26'd23451156;
ROM1[7186]<=26'd1954805; ROM2[7186]<=26'd11120995; ROM3[7186]<=26'd9746282; ROM4[7186]<=26'd23458799;
ROM1[7187]<=26'd1956575; ROM2[7187]<=26'd11124243; ROM3[7187]<=26'd9750938; ROM4[7187]<=26'd23463555;
ROM1[7188]<=26'd1956089; ROM2[7188]<=26'd11118961; ROM3[7188]<=26'd9745701; ROM4[7188]<=26'd23459661;
ROM1[7189]<=26'd1959737; ROM2[7189]<=26'd11115341; ROM3[7189]<=26'd9734889; ROM4[7189]<=26'd23454129;
ROM1[7190]<=26'd1969098; ROM2[7190]<=26'd11115419; ROM3[7190]<=26'd9730248; ROM4[7190]<=26'd23452864;
ROM1[7191]<=26'd1968658; ROM2[7191]<=26'd11115255; ROM3[7191]<=26'd9730848; ROM4[7191]<=26'd23453817;
ROM1[7192]<=26'd1960394; ROM2[7192]<=26'd11113720; ROM3[7192]<=26'd9732080; ROM4[7192]<=26'd23452470;
ROM1[7193]<=26'd1957302; ROM2[7193]<=26'd11115165; ROM3[7193]<=26'd9739955; ROM4[7193]<=26'd23456241;
ROM1[7194]<=26'd1959814; ROM2[7194]<=26'd11122525; ROM3[7194]<=26'd9749168; ROM4[7194]<=26'd23464260;
ROM1[7195]<=26'd1954645; ROM2[7195]<=26'd11121726; ROM3[7195]<=26'd9750449; ROM4[7195]<=26'd23463130;
ROM1[7196]<=26'd1952417; ROM2[7196]<=26'd11119546; ROM3[7196]<=26'd9747007; ROM4[7196]<=26'd23460595;
ROM1[7197]<=26'd1958973; ROM2[7197]<=26'd11119650; ROM3[7197]<=26'd9742092; ROM4[7197]<=26'd23458655;
ROM1[7198]<=26'd1963640; ROM2[7198]<=26'd11113480; ROM3[7198]<=26'd9730089; ROM4[7198]<=26'd23450558;
ROM1[7199]<=26'd1968697; ROM2[7199]<=26'd11116697; ROM3[7199]<=26'd9729781; ROM4[7199]<=26'd23451641;
ROM1[7200]<=26'd1968497; ROM2[7200]<=26'd11119485; ROM3[7200]<=26'd9734233; ROM4[7200]<=26'd23452605;
ROM1[7201]<=26'd1959575; ROM2[7201]<=26'd11118152; ROM3[7201]<=26'd9735492; ROM4[7201]<=26'd23452454;
ROM1[7202]<=26'd1957189; ROM2[7202]<=26'd11121404; ROM3[7202]<=26'd9741489; ROM4[7202]<=26'd23456728;
ROM1[7203]<=26'd1950340; ROM2[7203]<=26'd11118330; ROM3[7203]<=26'd9742665; ROM4[7203]<=26'd23454307;
ROM1[7204]<=26'd1951013; ROM2[7204]<=26'd11121113; ROM3[7204]<=26'd9746530; ROM4[7204]<=26'd23457701;
ROM1[7205]<=26'd1963489; ROM2[7205]<=26'd11125984; ROM3[7205]<=26'd9747066; ROM4[7205]<=26'd23460434;
ROM1[7206]<=26'd1974347; ROM2[7206]<=26'd11124175; ROM3[7206]<=26'd9738676; ROM4[7206]<=26'd23456550;
ROM1[7207]<=26'd1977410; ROM2[7207]<=26'd11120683; ROM3[7207]<=26'd9731530; ROM4[7207]<=26'd23454658;
ROM1[7208]<=26'd1970700; ROM2[7208]<=26'd11118900; ROM3[7208]<=26'd9729955; ROM4[7208]<=26'd23453822;
ROM1[7209]<=26'd1962709; ROM2[7209]<=26'd11116977; ROM3[7209]<=26'd9731900; ROM4[7209]<=26'd23453739;
ROM1[7210]<=26'd1954976; ROM2[7210]<=26'd11113319; ROM3[7210]<=26'd9732624; ROM4[7210]<=26'd23452954;
ROM1[7211]<=26'd1951205; ROM2[7211]<=26'd11115395; ROM3[7211]<=26'd9734588; ROM4[7211]<=26'd23454277;
ROM1[7212]<=26'd1953826; ROM2[7212]<=26'd11121502; ROM3[7212]<=26'd9740498; ROM4[7212]<=26'd23460264;
ROM1[7213]<=26'd1955927; ROM2[7213]<=26'd11122790; ROM3[7213]<=26'd9739257; ROM4[7213]<=26'd23460946;
ROM1[7214]<=26'd1962827; ROM2[7214]<=26'd11121741; ROM3[7214]<=26'd9731498; ROM4[7214]<=26'd23456675;
ROM1[7215]<=26'd1976923; ROM2[7215]<=26'd11125101; ROM3[7215]<=26'd9727899; ROM4[7215]<=26'd23458902;
ROM1[7216]<=26'd1977805; ROM2[7216]<=26'd11125492; ROM3[7216]<=26'd9728928; ROM4[7216]<=26'd23459827;
ROM1[7217]<=26'd1971151; ROM2[7217]<=26'd11123790; ROM3[7217]<=26'd9730988; ROM4[7217]<=26'd23459064;
ROM1[7218]<=26'd1964622; ROM2[7218]<=26'd11122683; ROM3[7218]<=26'd9732758; ROM4[7218]<=26'd23457939;
ROM1[7219]<=26'd1959102; ROM2[7219]<=26'd11122160; ROM3[7219]<=26'd9734248; ROM4[7219]<=26'd23456989;
ROM1[7220]<=26'd1960040; ROM2[7220]<=26'd11125735; ROM3[7220]<=26'd9740104; ROM4[7220]<=26'd23459552;
ROM1[7221]<=26'd1969625; ROM2[7221]<=26'd11131947; ROM3[7221]<=26'd9747200; ROM4[7221]<=26'd23465349;
ROM1[7222]<=26'd1981473; ROM2[7222]<=26'd11136563; ROM3[7222]<=26'd9748842; ROM4[7222]<=26'd23469773;
ROM1[7223]<=26'd1987626; ROM2[7223]<=26'd11132370; ROM3[7223]<=26'd9739545; ROM4[7223]<=26'd23464641;
ROM1[7224]<=26'd1983568; ROM2[7224]<=26'd11126390; ROM3[7224]<=26'd9731254; ROM4[7224]<=26'd23458646;
ROM1[7225]<=26'd1974506; ROM2[7225]<=26'd11123890; ROM3[7225]<=26'd9730537; ROM4[7225]<=26'd23455566;
ROM1[7226]<=26'd1968689; ROM2[7226]<=26'd11125139; ROM3[7226]<=26'd9734921; ROM4[7226]<=26'd23457568;
ROM1[7227]<=26'd1967831; ROM2[7227]<=26'd11128651; ROM3[7227]<=26'd9742915; ROM4[7227]<=26'd23462811;
ROM1[7228]<=26'd1955859; ROM2[7228]<=26'd11122292; ROM3[7228]<=26'd9739778; ROM4[7228]<=26'd23457344;
ROM1[7229]<=26'd1950591; ROM2[7229]<=26'd11119141; ROM3[7229]<=26'd9735551; ROM4[7229]<=26'd23452128;
ROM1[7230]<=26'd1954524; ROM2[7230]<=26'd11118695; ROM3[7230]<=26'd9731613; ROM4[7230]<=26'd23448470;
ROM1[7231]<=26'd1962208; ROM2[7231]<=26'd11117199; ROM3[7231]<=26'd9720987; ROM4[7231]<=26'd23443331;
ROM1[7232]<=26'd1973880; ROM2[7232]<=26'd11121503; ROM3[7232]<=26'd9719056; ROM4[7232]<=26'd23447183;
ROM1[7233]<=26'd1973570; ROM2[7233]<=26'd11121040; ROM3[7233]<=26'd9720895; ROM4[7233]<=26'd23449122;
ROM1[7234]<=26'd1969442; ROM2[7234]<=26'd11122475; ROM3[7234]<=26'd9726049; ROM4[7234]<=26'd23450963;
ROM1[7235]<=26'd1969890; ROM2[7235]<=26'd11127656; ROM3[7235]<=26'd9735762; ROM4[7235]<=26'd23457065;
ROM1[7236]<=26'd1964229; ROM2[7236]<=26'd11126836; ROM3[7236]<=26'd9737507; ROM4[7236]<=26'd23457056;
ROM1[7237]<=26'd1955322; ROM2[7237]<=26'd11122214; ROM3[7237]<=26'd9734137; ROM4[7237]<=26'd23452457;
ROM1[7238]<=26'd1953373; ROM2[7238]<=26'd11117630; ROM3[7238]<=26'd9728645; ROM4[7238]<=26'd23447790;
ROM1[7239]<=26'd1974223; ROM2[7239]<=26'd11127502; ROM3[7239]<=26'd9730910; ROM4[7239]<=26'd23455584;
ROM1[7240]<=26'd1993823; ROM2[7240]<=26'd11136469; ROM3[7240]<=26'd9736582; ROM4[7240]<=26'd23465846;
ROM1[7241]<=26'd1983339; ROM2[7241]<=26'd11126546; ROM3[7241]<=26'd9731243; ROM4[7241]<=26'd23459293;
ROM1[7242]<=26'd1976449; ROM2[7242]<=26'd11123847; ROM3[7242]<=26'd9733951; ROM4[7242]<=26'd23460738;
ROM1[7243]<=26'd1967737; ROM2[7243]<=26'd11121121; ROM3[7243]<=26'd9736338; ROM4[7243]<=26'd23461034;
ROM1[7244]<=26'd1958284; ROM2[7244]<=26'd11115975; ROM3[7244]<=26'd9734809; ROM4[7244]<=26'd23456400;
ROM1[7245]<=26'd1958781; ROM2[7245]<=26'd11122105; ROM3[7245]<=26'd9743544; ROM4[7245]<=26'd23462793;
ROM1[7246]<=26'd1962118; ROM2[7246]<=26'd11127158; ROM3[7246]<=26'd9749881; ROM4[7246]<=26'd23468274;
ROM1[7247]<=26'd1964181; ROM2[7247]<=26'd11121111; ROM3[7247]<=26'd9741492; ROM4[7247]<=26'd23462897;
ROM1[7248]<=26'd1970138; ROM2[7248]<=26'd11115971; ROM3[7248]<=26'd9729567; ROM4[7248]<=26'd23456059;
ROM1[7249]<=26'd1981870; ROM2[7249]<=26'd11122936; ROM3[7249]<=26'd9734620; ROM4[7249]<=26'd23462952;
ROM1[7250]<=26'd1982633; ROM2[7250]<=26'd11127108; ROM3[7250]<=26'd9740802; ROM4[7250]<=26'd23467632;
ROM1[7251]<=26'd1971904; ROM2[7251]<=26'd11124103; ROM3[7251]<=26'd9742548; ROM4[7251]<=26'd23465528;
ROM1[7252]<=26'd1961369; ROM2[7252]<=26'd11120945; ROM3[7252]<=26'd9741248; ROM4[7252]<=26'd23462390;
ROM1[7253]<=26'd1954515; ROM2[7253]<=26'd11119650; ROM3[7253]<=26'd9740423; ROM4[7253]<=26'd23458910;
ROM1[7254]<=26'd1951914; ROM2[7254]<=26'd11117259; ROM3[7254]<=26'd9737554; ROM4[7254]<=26'd23455667;
ROM1[7255]<=26'd1959155; ROM2[7255]<=26'd11119598; ROM3[7255]<=26'd9737300; ROM4[7255]<=26'd23456054;
ROM1[7256]<=26'd1976776; ROM2[7256]<=26'd11125282; ROM3[7256]<=26'd9737151; ROM4[7256]<=26'd23459553;
ROM1[7257]<=26'd1983034; ROM2[7257]<=26'd11125223; ROM3[7257]<=26'd9731540; ROM4[7257]<=26'd23458987;
ROM1[7258]<=26'd1975414; ROM2[7258]<=26'd11120740; ROM3[7258]<=26'd9729362; ROM4[7258]<=26'd23455830;
ROM1[7259]<=26'd1966877; ROM2[7259]<=26'd11118427; ROM3[7259]<=26'd9732889; ROM4[7259]<=26'd23453995;
ROM1[7260]<=26'd1965850; ROM2[7260]<=26'd11122092; ROM3[7260]<=26'd9742180; ROM4[7260]<=26'd23457544;
ROM1[7261]<=26'd1961033; ROM2[7261]<=26'd11122066; ROM3[7261]<=26'd9745677; ROM4[7261]<=26'd23459353;
ROM1[7262]<=26'd1955389; ROM2[7262]<=26'd11118274; ROM3[7262]<=26'd9744890; ROM4[7262]<=26'd23456110;
ROM1[7263]<=26'd1961250; ROM2[7263]<=26'd11121241; ROM3[7263]<=26'd9745653; ROM4[7263]<=26'd23458841;
ROM1[7264]<=26'd1973447; ROM2[7264]<=26'd11125226; ROM3[7264]<=26'd9743834; ROM4[7264]<=26'd23461369;
ROM1[7265]<=26'd1987418; ROM2[7265]<=26'd11128992; ROM3[7265]<=26'd9743394; ROM4[7265]<=26'd23463730;
ROM1[7266]<=26'd1987515; ROM2[7266]<=26'd11130665; ROM3[7266]<=26'd9745052; ROM4[7266]<=26'd23466923;
ROM1[7267]<=26'd1978310; ROM2[7267]<=26'd11126238; ROM3[7267]<=26'd9744687; ROM4[7267]<=26'd23465833;
ROM1[7268]<=26'd1974356; ROM2[7268]<=26'd11127026; ROM3[7268]<=26'd9750571; ROM4[7268]<=26'd23469902;
ROM1[7269]<=26'd1976490; ROM2[7269]<=26'd11132491; ROM3[7269]<=26'd9756783; ROM4[7269]<=26'd23476179;
ROM1[7270]<=26'd1973432; ROM2[7270]<=26'd11133619; ROM3[7270]<=26'd9756174; ROM4[7270]<=26'd23476221;
ROM1[7271]<=26'd1977205; ROM2[7271]<=26'd11136754; ROM3[7271]<=26'd9757688; ROM4[7271]<=26'd23479390;
ROM1[7272]<=26'd1983269; ROM2[7272]<=26'd11134888; ROM3[7272]<=26'd9751498; ROM4[7272]<=26'd23476595;
ROM1[7273]<=26'd1986243; ROM2[7273]<=26'd11126256; ROM3[7273]<=26'd9736699; ROM4[7273]<=26'd23467181;
ROM1[7274]<=26'd1986155; ROM2[7274]<=26'd11123013; ROM3[7274]<=26'd9732453; ROM4[7274]<=26'd23462830;
ROM1[7275]<=26'd1983350; ROM2[7275]<=26'd11126915; ROM3[7275]<=26'd9737335; ROM4[7275]<=26'd23464349;
ROM1[7276]<=26'd1976762; ROM2[7276]<=26'd11129584; ROM3[7276]<=26'd9743593; ROM4[7276]<=26'd23466453;
ROM1[7277]<=26'd1965007; ROM2[7277]<=26'd11124399; ROM3[7277]<=26'd9741303; ROM4[7277]<=26'd23461528;
ROM1[7278]<=26'd1961027; ROM2[7278]<=26'd11125332; ROM3[7278]<=26'd9742444; ROM4[7278]<=26'd23461045;
ROM1[7279]<=26'd1957145; ROM2[7279]<=26'd11122410; ROM3[7279]<=26'd9739406; ROM4[7279]<=26'd23458144;
ROM1[7280]<=26'd1956572; ROM2[7280]<=26'd11115063; ROM3[7280]<=26'd9729439; ROM4[7280]<=26'd23451224;
ROM1[7281]<=26'd1973258; ROM2[7281]<=26'd11121125; ROM3[7281]<=26'd9730426; ROM4[7281]<=26'd23454953;
ROM1[7282]<=26'd1988298; ROM2[7282]<=26'd11129613; ROM3[7282]<=26'd9737200; ROM4[7282]<=26'd23463204;
ROM1[7283]<=26'd1986428; ROM2[7283]<=26'd11129119; ROM3[7283]<=26'd9738401; ROM4[7283]<=26'd23462976;
ROM1[7284]<=26'd1976212; ROM2[7284]<=26'd11124027; ROM3[7284]<=26'd9736951; ROM4[7284]<=26'd23458870;
ROM1[7285]<=26'd1970250; ROM2[7285]<=26'd11122978; ROM3[7285]<=26'd9741219; ROM4[7285]<=26'd23460685;
ROM1[7286]<=26'd1962728; ROM2[7286]<=26'd11119854; ROM3[7286]<=26'd9740940; ROM4[7286]<=26'd23459467;
ROM1[7287]<=26'd1958882; ROM2[7287]<=26'd11118846; ROM3[7287]<=26'd9740943; ROM4[7287]<=26'd23458438;
ROM1[7288]<=26'd1966303; ROM2[7288]<=26'd11123406; ROM3[7288]<=26'd9744214; ROM4[7288]<=26'd23462245;
ROM1[7289]<=26'd1979212; ROM2[7289]<=26'd11127557; ROM3[7289]<=26'd9743694; ROM4[7289]<=26'd23464292;
ROM1[7290]<=26'd1985596; ROM2[7290]<=26'd11125396; ROM3[7290]<=26'd9736403; ROM4[7290]<=26'd23460389;
ROM1[7291]<=26'd1980680; ROM2[7291]<=26'd11121429; ROM3[7291]<=26'd9734455; ROM4[7291]<=26'd23458813;
ROM1[7292]<=26'd1979494; ROM2[7292]<=26'd11125792; ROM3[7292]<=26'd9742717; ROM4[7292]<=26'd23464730;
ROM1[7293]<=26'd1975653; ROM2[7293]<=26'd11128630; ROM3[7293]<=26'd9747499; ROM4[7293]<=26'd23467019;
ROM1[7294]<=26'd1970227; ROM2[7294]<=26'd11128195; ROM3[7294]<=26'd9748076; ROM4[7294]<=26'd23467037;
ROM1[7295]<=26'd1964717; ROM2[7295]<=26'd11128178; ROM3[7295]<=26'd9749766; ROM4[7295]<=26'd23467367;
ROM1[7296]<=26'd1962367; ROM2[7296]<=26'd11124645; ROM3[7296]<=26'd9747668; ROM4[7296]<=26'd23464424;
ROM1[7297]<=26'd1969028; ROM2[7297]<=26'd11122975; ROM3[7297]<=26'd9742188; ROM4[7297]<=26'd23462853;
ROM1[7298]<=26'd1985371; ROM2[7298]<=26'd11127786; ROM3[7298]<=26'd9741808; ROM4[7298]<=26'd23467045;
ROM1[7299]<=26'd1992254; ROM2[7299]<=26'd11131537; ROM3[7299]<=26'd9745868; ROM4[7299]<=26'd23469963;
ROM1[7300]<=26'd1985397; ROM2[7300]<=26'd11131046; ROM3[7300]<=26'd9745557; ROM4[7300]<=26'd23469480;
ROM1[7301]<=26'd1974730; ROM2[7301]<=26'd11123595; ROM3[7301]<=26'd9744833; ROM4[7301]<=26'd23466410;
ROM1[7302]<=26'd1964003; ROM2[7302]<=26'd11114880; ROM3[7302]<=26'd9743780; ROM4[7302]<=26'd23461609;
ROM1[7303]<=26'd1953781; ROM2[7303]<=26'd11108266; ROM3[7303]<=26'd9741508; ROM4[7303]<=26'd23457101;
ROM1[7304]<=26'd1954194; ROM2[7304]<=26'd11111282; ROM3[7304]<=26'd9744798; ROM4[7304]<=26'd23459142;
ROM1[7305]<=26'd1966050; ROM2[7305]<=26'd11118649; ROM3[7305]<=26'd9748397; ROM4[7305]<=26'd23464416;
ROM1[7306]<=26'd1976664; ROM2[7306]<=26'd11117108; ROM3[7306]<=26'd9742675; ROM4[7306]<=26'd23462160;
ROM1[7307]<=26'd1983516; ROM2[7307]<=26'd11119135; ROM3[7307]<=26'd9739551; ROM4[7307]<=26'd23461621;
ROM1[7308]<=26'd1987360; ROM2[7308]<=26'd11126085; ROM3[7308]<=26'd9747461; ROM4[7308]<=26'd23468835;
ROM1[7309]<=26'd1978013; ROM2[7309]<=26'd11124242; ROM3[7309]<=26'd9749076; ROM4[7309]<=26'd23468045;
ROM1[7310]<=26'd1964771; ROM2[7310]<=26'd11117418; ROM3[7310]<=26'd9745211; ROM4[7310]<=26'd23461482;
ROM1[7311]<=26'd1959936; ROM2[7311]<=26'd11117670; ROM3[7311]<=26'd9748390; ROM4[7311]<=26'd23463387;
ROM1[7312]<=26'd1954782; ROM2[7312]<=26'd11116872; ROM3[7312]<=26'd9747181; ROM4[7312]<=26'd23461858;
ROM1[7313]<=26'd1960180; ROM2[7313]<=26'd11118270; ROM3[7313]<=26'd9748190; ROM4[7313]<=26'd23462429;
ROM1[7314]<=26'd1978074; ROM2[7314]<=26'd11126737; ROM3[7314]<=26'd9751523; ROM4[7314]<=26'd23468995;
ROM1[7315]<=26'd1987859; ROM2[7315]<=26'd11125883; ROM3[7315]<=26'd9744012; ROM4[7315]<=26'd23467510;
ROM1[7316]<=26'd1987117; ROM2[7316]<=26'd11122980; ROM3[7316]<=26'd9743105; ROM4[7316]<=26'd23466222;
ROM1[7317]<=26'd1982051; ROM2[7317]<=26'd11126633; ROM3[7317]<=26'd9746621; ROM4[7317]<=26'd23467047;
ROM1[7318]<=26'd1971761; ROM2[7318]<=26'd11121520; ROM3[7318]<=26'd9742988; ROM4[7318]<=26'd23463208;
ROM1[7319]<=26'd1968512; ROM2[7319]<=26'd11120151; ROM3[7319]<=26'd9747072; ROM4[7319]<=26'd23464147;
ROM1[7320]<=26'd1959870; ROM2[7320]<=26'd11116820; ROM3[7320]<=26'd9747902; ROM4[7320]<=26'd23462383;
ROM1[7321]<=26'd1954386; ROM2[7321]<=26'd11112185; ROM3[7321]<=26'd9741644; ROM4[7321]<=26'd23458642;
ROM1[7322]<=26'd1967304; ROM2[7322]<=26'd11119201; ROM3[7322]<=26'd9742660; ROM4[7322]<=26'd23461727;
ROM1[7323]<=26'd1981188; ROM2[7323]<=26'd11121849; ROM3[7323]<=26'd9738999; ROM4[7323]<=26'd23462793;
ROM1[7324]<=26'd1983384; ROM2[7324]<=26'd11120837; ROM3[7324]<=26'd9734702; ROM4[7324]<=26'd23461121;
ROM1[7325]<=26'd1983302; ROM2[7325]<=26'd11125056; ROM3[7325]<=26'd9741630; ROM4[7325]<=26'd23466280;
ROM1[7326]<=26'd1978639; ROM2[7326]<=26'd11127876; ROM3[7326]<=26'd9750431; ROM4[7326]<=26'd23472318;
ROM1[7327]<=26'd1967734; ROM2[7327]<=26'd11122771; ROM3[7327]<=26'd9746532; ROM4[7327]<=26'd23467114;
ROM1[7328]<=26'd1958539; ROM2[7328]<=26'd11119874; ROM3[7328]<=26'd9743343; ROM4[7328]<=26'd23462516;
ROM1[7329]<=26'd1951955; ROM2[7329]<=26'd11113377; ROM3[7329]<=26'd9739861; ROM4[7329]<=26'd23457527;
ROM1[7330]<=26'd1954969; ROM2[7330]<=26'd11110822; ROM3[7330]<=26'd9735637; ROM4[7330]<=26'd23456186;
ROM1[7331]<=26'd1969600; ROM2[7331]<=26'd11116791; ROM3[7331]<=26'd9734865; ROM4[7331]<=26'd23460200;
ROM1[7332]<=26'd1981841; ROM2[7332]<=26'd11121269; ROM3[7332]<=26'd9738862; ROM4[7332]<=26'd23465252;
ROM1[7333]<=26'd1980255; ROM2[7333]<=26'd11122559; ROM3[7333]<=26'd9740107; ROM4[7333]<=26'd23466616;
ROM1[7334]<=26'd1966050; ROM2[7334]<=26'd11114815; ROM3[7334]<=26'd9733787; ROM4[7334]<=26'd23458805;
ROM1[7335]<=26'd1957261; ROM2[7335]<=26'd11111366; ROM3[7335]<=26'd9732372; ROM4[7335]<=26'd23454661;
ROM1[7336]<=26'd1954993; ROM2[7336]<=26'd11112559; ROM3[7336]<=26'd9734024; ROM4[7336]<=26'd23454958;
ROM1[7337]<=26'd1956076; ROM2[7337]<=26'd11115740; ROM3[7337]<=26'd9739777; ROM4[7337]<=26'd23458747;
ROM1[7338]<=26'd1963804; ROM2[7338]<=26'd11120643; ROM3[7338]<=26'd9742404; ROM4[7338]<=26'd23462434;
ROM1[7339]<=26'd1972200; ROM2[7339]<=26'd11118957; ROM3[7339]<=26'd9733893; ROM4[7339]<=26'd23459214;
ROM1[7340]<=26'd1978121; ROM2[7340]<=26'd11114757; ROM3[7340]<=26'd9726775; ROM4[7340]<=26'd23455647;
ROM1[7341]<=26'd1974743; ROM2[7341]<=26'd11113298; ROM3[7341]<=26'd9724832; ROM4[7341]<=26'd23453179;
ROM1[7342]<=26'd1971312; ROM2[7342]<=26'd11118265; ROM3[7342]<=26'd9728357; ROM4[7342]<=26'd23454967;
ROM1[7343]<=26'd1965280; ROM2[7343]<=26'd11119398; ROM3[7343]<=26'd9733690; ROM4[7343]<=26'd23456677;
ROM1[7344]<=26'd1957225; ROM2[7344]<=26'd11117625; ROM3[7344]<=26'd9735038; ROM4[7344]<=26'd23456765;
ROM1[7345]<=26'd1956211; ROM2[7345]<=26'd11120237; ROM3[7345]<=26'd9739640; ROM4[7345]<=26'd23460077;
ROM1[7346]<=26'd1958351; ROM2[7346]<=26'd11119877; ROM3[7346]<=26'd9740780; ROM4[7346]<=26'd23460409;
ROM1[7347]<=26'd1965587; ROM2[7347]<=26'd11119011; ROM3[7347]<=26'd9737194; ROM4[7347]<=26'd23458297;
ROM1[7348]<=26'd1972126; ROM2[7348]<=26'd11113815; ROM3[7348]<=26'd9725547; ROM4[7348]<=26'd23450857;
ROM1[7349]<=26'd1970207; ROM2[7349]<=26'd11110165; ROM3[7349]<=26'd9720399; ROM4[7349]<=26'd23446920;
ROM1[7350]<=26'd1966398; ROM2[7350]<=26'd11111042; ROM3[7350]<=26'd9725621; ROM4[7350]<=26'd23450508;
ROM1[7351]<=26'd1962411; ROM2[7351]<=26'd11112597; ROM3[7351]<=26'd9731426; ROM4[7351]<=26'd23454235;
ROM1[7352]<=26'd1960307; ROM2[7352]<=26'd11117895; ROM3[7352]<=26'd9737960; ROM4[7352]<=26'd23458224;
ROM1[7353]<=26'd1954450; ROM2[7353]<=26'd11116359; ROM3[7353]<=26'd9741507; ROM4[7353]<=26'd23458356;
ROM1[7354]<=26'd1954471; ROM2[7354]<=26'd11118675; ROM3[7354]<=26'd9745205; ROM4[7354]<=26'd23462331;
ROM1[7355]<=26'd1959884; ROM2[7355]<=26'd11119677; ROM3[7355]<=26'd9743071; ROM4[7355]<=26'd23463491;
ROM1[7356]<=26'd1973691; ROM2[7356]<=26'd11119871; ROM3[7356]<=26'd9736289; ROM4[7356]<=26'd23462171;
ROM1[7357]<=26'd1982859; ROM2[7357]<=26'd11124720; ROM3[7357]<=26'd9734544; ROM4[7357]<=26'd23464908;
ROM1[7358]<=26'd1980472; ROM2[7358]<=26'd11126566; ROM3[7358]<=26'd9738578; ROM4[7358]<=26'd23465917;
ROM1[7359]<=26'd1975443; ROM2[7359]<=26'd11126410; ROM3[7359]<=26'd9741999; ROM4[7359]<=26'd23465277;
ROM1[7360]<=26'd1969197; ROM2[7360]<=26'd11124946; ROM3[7360]<=26'd9744496; ROM4[7360]<=26'd23466461;
ROM1[7361]<=26'd1961530; ROM2[7361]<=26'd11122502; ROM3[7361]<=26'd9744222; ROM4[7361]<=26'd23464446;
ROM1[7362]<=26'd1953578; ROM2[7362]<=26'd11118862; ROM3[7362]<=26'd9739431; ROM4[7362]<=26'd23459783;
ROM1[7363]<=26'd1957928; ROM2[7363]<=26'd11121158; ROM3[7363]<=26'd9738793; ROM4[7363]<=26'd23461282;
ROM1[7364]<=26'd1972959; ROM2[7364]<=26'd11126011; ROM3[7364]<=26'd9739545; ROM4[7364]<=26'd23464050;
ROM1[7365]<=26'd1983271; ROM2[7365]<=26'd11125234; ROM3[7365]<=26'd9734468; ROM4[7365]<=26'd23462413;
ROM1[7366]<=26'd1981116; ROM2[7366]<=26'd11123110; ROM3[7366]<=26'd9731500; ROM4[7366]<=26'd23460386;
ROM1[7367]<=26'd1976403; ROM2[7367]<=26'd11124217; ROM3[7367]<=26'd9736075; ROM4[7367]<=26'd23463357;
ROM1[7368]<=26'd1970653; ROM2[7368]<=26'd11124481; ROM3[7368]<=26'd9741083; ROM4[7368]<=26'd23465452;
ROM1[7369]<=26'd1969453; ROM2[7369]<=26'd11126211; ROM3[7369]<=26'd9745419; ROM4[7369]<=26'd23467835;
ROM1[7370]<=26'd1966880; ROM2[7370]<=26'd11127179; ROM3[7370]<=26'd9747573; ROM4[7370]<=26'd23468560;
ROM1[7371]<=26'd1965924; ROM2[7371]<=26'd11124833; ROM3[7371]<=26'd9746454; ROM4[7371]<=26'd23465576;
ROM1[7372]<=26'd1975886; ROM2[7372]<=26'd11127493; ROM3[7372]<=26'd9744239; ROM4[7372]<=26'd23465416;
ROM1[7373]<=26'd1989367; ROM2[7373]<=26'd11128903; ROM3[7373]<=26'd9737921; ROM4[7373]<=26'd23465526;
ROM1[7374]<=26'd1992858; ROM2[7374]<=26'd11130723; ROM3[7374]<=26'd9737978; ROM4[7374]<=26'd23466384;
ROM1[7375]<=26'd1985997; ROM2[7375]<=26'd11130625; ROM3[7375]<=26'd9739756; ROM4[7375]<=26'd23468072;
ROM1[7376]<=26'd1972268; ROM2[7376]<=26'd11124391; ROM3[7376]<=26'd9737761; ROM4[7376]<=26'd23464641;
ROM1[7377]<=26'd1963478; ROM2[7377]<=26'd11122124; ROM3[7377]<=26'd9739902; ROM4[7377]<=26'd23462059;
ROM1[7378]<=26'd1958665; ROM2[7378]<=26'd11123018; ROM3[7378]<=26'd9744137; ROM4[7378]<=26'd23463973;
ROM1[7379]<=26'd1956649; ROM2[7379]<=26'd11123147; ROM3[7379]<=26'd9741820; ROM4[7379]<=26'd23461645;
ROM1[7380]<=26'd1956951; ROM2[7380]<=26'd11118082; ROM3[7380]<=26'd9731821; ROM4[7380]<=26'd23455261;
ROM1[7381]<=26'd1966843; ROM2[7381]<=26'd11117113; ROM3[7381]<=26'd9725268; ROM4[7381]<=26'd23454603;
ROM1[7382]<=26'd1975710; ROM2[7382]<=26'd11116759; ROM3[7382]<=26'd9722562; ROM4[7382]<=26'd23454690;
ROM1[7383]<=26'd1973521; ROM2[7383]<=26'd11117120; ROM3[7383]<=26'd9725004; ROM4[7383]<=26'd23455566;
ROM1[7384]<=26'd1965358; ROM2[7384]<=26'd11116673; ROM3[7384]<=26'd9728186; ROM4[7384]<=26'd23454371;
ROM1[7385]<=26'd1955225; ROM2[7385]<=26'd11113738; ROM3[7385]<=26'd9727917; ROM4[7385]<=26'd23452224;
ROM1[7386]<=26'd1953772; ROM2[7386]<=26'd11116546; ROM3[7386]<=26'd9733238; ROM4[7386]<=26'd23456195;
ROM1[7387]<=26'd1954983; ROM2[7387]<=26'd11119317; ROM3[7387]<=26'd9740407; ROM4[7387]<=26'd23459800;
ROM1[7388]<=26'd1959087; ROM2[7388]<=26'd11121349; ROM3[7388]<=26'd9740020; ROM4[7388]<=26'd23460629;
ROM1[7389]<=26'd1961700; ROM2[7389]<=26'd11111698; ROM3[7389]<=26'd9725030; ROM4[7389]<=26'd23451514;
ROM1[7390]<=26'd1966490; ROM2[7390]<=26'd11106492; ROM3[7390]<=26'd9713576; ROM4[7390]<=26'd23444264;
ROM1[7391]<=26'd1966261; ROM2[7391]<=26'd11109763; ROM3[7391]<=26'd9713395; ROM4[7391]<=26'd23444464;
ROM1[7392]<=26'd1964604; ROM2[7392]<=26'd11113728; ROM3[7392]<=26'd9720291; ROM4[7392]<=26'd23449706;
ROM1[7393]<=26'd1967288; ROM2[7393]<=26'd11123198; ROM3[7393]<=26'd9732601; ROM4[7393]<=26'd23457877;
ROM1[7394]<=26'd1960293; ROM2[7394]<=26'd11122663; ROM3[7394]<=26'd9734631; ROM4[7394]<=26'd23458960;
ROM1[7395]<=26'd1953568; ROM2[7395]<=26'd11119116; ROM3[7395]<=26'd9735623; ROM4[7395]<=26'd23458801;
ROM1[7396]<=26'd1961815; ROM2[7396]<=26'd11126495; ROM3[7396]<=26'd9739505; ROM4[7396]<=26'd23464003;
ROM1[7397]<=26'd1972924; ROM2[7397]<=26'd11129203; ROM3[7397]<=26'd9735186; ROM4[7397]<=26'd23464523;
ROM1[7398]<=26'd1979248; ROM2[7398]<=26'd11124345; ROM3[7398]<=26'd9726675; ROM4[7398]<=26'd23459751;
ROM1[7399]<=26'd1981922; ROM2[7399]<=26'd11123150; ROM3[7399]<=26'd9723878; ROM4[7399]<=26'd23459179;
ROM1[7400]<=26'd1976537; ROM2[7400]<=26'd11120375; ROM3[7400]<=26'd9724916; ROM4[7400]<=26'd23458661;
ROM1[7401]<=26'd1971698; ROM2[7401]<=26'd11121375; ROM3[7401]<=26'd9730711; ROM4[7401]<=26'd23461376;
ROM1[7402]<=26'd1971935; ROM2[7402]<=26'd11125434; ROM3[7402]<=26'd9739192; ROM4[7402]<=26'd23466991;
ROM1[7403]<=26'd1964161; ROM2[7403]<=26'd11123906; ROM3[7403]<=26'd9740679; ROM4[7403]<=26'd23465925;
ROM1[7404]<=26'd1961838; ROM2[7404]<=26'd11122005; ROM3[7404]<=26'd9741599; ROM4[7404]<=26'd23465920;
ROM1[7405]<=26'd1968574; ROM2[7405]<=26'd11124281; ROM3[7405]<=26'd9741314; ROM4[7405]<=26'd23466968;
ROM1[7406]<=26'd1977835; ROM2[7406]<=26'd11122232; ROM3[7406]<=26'd9732248; ROM4[7406]<=26'd23459706;
ROM1[7407]<=26'd1980492; ROM2[7407]<=26'd11117797; ROM3[7407]<=26'd9725990; ROM4[7407]<=26'd23456248;
ROM1[7408]<=26'd1979325; ROM2[7408]<=26'd11120937; ROM3[7408]<=26'd9730898; ROM4[7408]<=26'd23461195;
ROM1[7409]<=26'd1975161; ROM2[7409]<=26'd11122575; ROM3[7409]<=26'd9737912; ROM4[7409]<=26'd23464141;
ROM1[7410]<=26'd1969835; ROM2[7410]<=26'd11122142; ROM3[7410]<=26'd9743078; ROM4[7410]<=26'd23467445;
ROM1[7411]<=26'd1969795; ROM2[7411]<=26'd11127462; ROM3[7411]<=26'd9754258; ROM4[7411]<=26'd23473718;
ROM1[7412]<=26'd1972197; ROM2[7412]<=26'd11133182; ROM3[7412]<=26'd9763566; ROM4[7412]<=26'd23481456;
ROM1[7413]<=26'd1972136; ROM2[7413]<=26'd11131963; ROM3[7413]<=26'd9759939; ROM4[7413]<=26'd23480775;
ROM1[7414]<=26'd1979804; ROM2[7414]<=26'd11130441; ROM3[7414]<=26'd9751789; ROM4[7414]<=26'd23475789;
ROM1[7415]<=26'd1991945; ROM2[7415]<=26'd11131576; ROM3[7415]<=26'd9744683; ROM4[7415]<=26'd23474237;
ROM1[7416]<=26'd1988615; ROM2[7416]<=26'd11130701; ROM3[7416]<=26'd9741123; ROM4[7416]<=26'd23470533;
ROM1[7417]<=26'd1984649; ROM2[7417]<=26'd11133728; ROM3[7417]<=26'd9749000; ROM4[7417]<=26'd23473278;
ROM1[7418]<=26'd1979834; ROM2[7418]<=26'd11135146; ROM3[7418]<=26'd9753734; ROM4[7418]<=26'd23476204;
ROM1[7419]<=26'd1968304; ROM2[7419]<=26'd11129445; ROM3[7419]<=26'd9748645; ROM4[7419]<=26'd23470541;
ROM1[7420]<=26'd1959451; ROM2[7420]<=26'd11123961; ROM3[7420]<=26'd9745077; ROM4[7420]<=26'd23464541;
ROM1[7421]<=26'd1959804; ROM2[7421]<=26'd11121792; ROM3[7421]<=26'd9741708; ROM4[7421]<=26'd23461136;
ROM1[7422]<=26'd1969304; ROM2[7422]<=26'd11125342; ROM3[7422]<=26'd9738626; ROM4[7422]<=26'd23460904;
ROM1[7423]<=26'd1983898; ROM2[7423]<=26'd11128363; ROM3[7423]<=26'd9735035; ROM4[7423]<=26'd23462846;
ROM1[7424]<=26'd1985609; ROM2[7424]<=26'd11126747; ROM3[7424]<=26'd9731908; ROM4[7424]<=26'd23462389;
ROM1[7425]<=26'd1978345; ROM2[7425]<=26'd11123669; ROM3[7425]<=26'd9730509; ROM4[7425]<=26'd23460072;
ROM1[7426]<=26'd1970506; ROM2[7426]<=26'd11122278; ROM3[7426]<=26'd9731946; ROM4[7426]<=26'd23460082;
ROM1[7427]<=26'd1967623; ROM2[7427]<=26'd11123732; ROM3[7427]<=26'd9735591; ROM4[7427]<=26'd23461446;
ROM1[7428]<=26'd1961953; ROM2[7428]<=26'd11122912; ROM3[7428]<=26'd9735199; ROM4[7428]<=26'd23458053;
ROM1[7429]<=26'd1960926; ROM2[7429]<=26'd11124742; ROM3[7429]<=26'd9734936; ROM4[7429]<=26'd23458245;
ROM1[7430]<=26'd1968493; ROM2[7430]<=26'd11126263; ROM3[7430]<=26'd9732951; ROM4[7430]<=26'd23458160;
ROM1[7431]<=26'd1979006; ROM2[7431]<=26'd11125743; ROM3[7431]<=26'd9722981; ROM4[7431]<=26'd23454191;
ROM1[7432]<=26'd1988640; ROM2[7432]<=26'd11130420; ROM3[7432]<=26'd9722493; ROM4[7432]<=26'd23457435;
ROM1[7433]<=26'd1987375; ROM2[7433]<=26'd11134422; ROM3[7433]<=26'd9726172; ROM4[7433]<=26'd23460073;
ROM1[7434]<=26'd1979631; ROM2[7434]<=26'd11133392; ROM3[7434]<=26'd9727165; ROM4[7434]<=26'd23460099;
ROM1[7435]<=26'd1968278; ROM2[7435]<=26'd11127916; ROM3[7435]<=26'd9724641; ROM4[7435]<=26'd23455104;
ROM1[7436]<=26'd1952709; ROM2[7436]<=26'd11120059; ROM3[7436]<=26'd9719931; ROM4[7436]<=26'd23447678;
ROM1[7437]<=26'd1947130; ROM2[7437]<=26'd11117529; ROM3[7437]<=26'd9719237; ROM4[7437]<=26'd23444995;
ROM1[7438]<=26'd1954634; ROM2[7438]<=26'd11120649; ROM3[7438]<=26'd9719584; ROM4[7438]<=26'd23445489;
ROM1[7439]<=26'd1968102; ROM2[7439]<=26'd11122962; ROM3[7439]<=26'd9716970; ROM4[7439]<=26'd23447535;
ROM1[7440]<=26'd1981018; ROM2[7440]<=26'd11122667; ROM3[7440]<=26'd9714603; ROM4[7440]<=26'd23447532;
ROM1[7441]<=26'd1984152; ROM2[7441]<=26'd11124342; ROM3[7441]<=26'd9718592; ROM4[7441]<=26'd23451650;
ROM1[7442]<=26'd1979970; ROM2[7442]<=26'd11126114; ROM3[7442]<=26'd9725151; ROM4[7442]<=26'd23454962;
ROM1[7443]<=26'd1977517; ROM2[7443]<=26'd11130200; ROM3[7443]<=26'd9736684; ROM4[7443]<=26'd23459832;
ROM1[7444]<=26'd1972188; ROM2[7444]<=26'd11131117; ROM3[7444]<=26'd9738992; ROM4[7444]<=26'd23462158;
ROM1[7445]<=26'd1955396; ROM2[7445]<=26'd11118993; ROM3[7445]<=26'd9729436; ROM4[7445]<=26'd23451534;
ROM1[7446]<=26'd1950752; ROM2[7446]<=26'd11114171; ROM3[7446]<=26'd9726054; ROM4[7446]<=26'd23447152;
ROM1[7447]<=26'd1960890; ROM2[7447]<=26'd11117197; ROM3[7447]<=26'd9725391; ROM4[7447]<=26'd23450486;
ROM1[7448]<=26'd1973965; ROM2[7448]<=26'd11118979; ROM3[7448]<=26'd9721102; ROM4[7448]<=26'd23451589;
ROM1[7449]<=26'd1981781; ROM2[7449]<=26'd11124014; ROM3[7449]<=26'd9725117; ROM4[7449]<=26'd23456632;
ROM1[7450]<=26'd1984046; ROM2[7450]<=26'd11132198; ROM3[7450]<=26'd9736172; ROM4[7450]<=26'd23465600;
ROM1[7451]<=26'd1977037; ROM2[7451]<=26'd11132754; ROM3[7451]<=26'd9739597; ROM4[7451]<=26'd23465965;
ROM1[7452]<=26'd1971062; ROM2[7452]<=26'd11131218; ROM3[7452]<=26'd9741398; ROM4[7452]<=26'd23465319;
ROM1[7453]<=26'd1967091; ROM2[7453]<=26'd11131412; ROM3[7453]<=26'd9745673; ROM4[7453]<=26'd23466997;
ROM1[7454]<=26'd1961990; ROM2[7454]<=26'd11128154; ROM3[7454]<=26'd9741737; ROM4[7454]<=26'd23464077;
ROM1[7455]<=26'd1967241; ROM2[7455]<=26'd11126633; ROM3[7455]<=26'd9738578; ROM4[7455]<=26'd23464926;
ROM1[7456]<=26'd1980396; ROM2[7456]<=26'd11126646; ROM3[7456]<=26'd9735679; ROM4[7456]<=26'd23464871;
ROM1[7457]<=26'd1986022; ROM2[7457]<=26'd11128629; ROM3[7457]<=26'd9732428; ROM4[7457]<=26'd23465093;
ROM1[7458]<=26'd1982743; ROM2[7458]<=26'd11128953; ROM3[7458]<=26'd9735079; ROM4[7458]<=26'd23465969;
ROM1[7459]<=26'd1974804; ROM2[7459]<=26'd11126038; ROM3[7459]<=26'd9737867; ROM4[7459]<=26'd23463983;
ROM1[7460]<=26'd1968875; ROM2[7460]<=26'd11126284; ROM3[7460]<=26'd9741016; ROM4[7460]<=26'd23465353;
ROM1[7461]<=26'd1963429; ROM2[7461]<=26'd11124942; ROM3[7461]<=26'd9742702; ROM4[7461]<=26'd23464226;
ROM1[7462]<=26'd1957801; ROM2[7462]<=26'd11122815; ROM3[7462]<=26'd9742742; ROM4[7462]<=26'd23462565;
ROM1[7463]<=26'd1960840; ROM2[7463]<=26'd11123599; ROM3[7463]<=26'd9742429; ROM4[7463]<=26'd23461562;
ROM1[7464]<=26'd1975426; ROM2[7464]<=26'd11127837; ROM3[7464]<=26'd9740110; ROM4[7464]<=26'd23462029;
ROM1[7465]<=26'd1986833; ROM2[7465]<=26'd11130951; ROM3[7465]<=26'd9736391; ROM4[7465]<=26'd23463149;
ROM1[7466]<=26'd1983997; ROM2[7466]<=26'd11128443; ROM3[7466]<=26'd9734622; ROM4[7466]<=26'd23460357;
ROM1[7467]<=26'd1977343; ROM2[7467]<=26'd11128201; ROM3[7467]<=26'd9736604; ROM4[7467]<=26'd23459723;
ROM1[7468]<=26'd1967904; ROM2[7468]<=26'd11125253; ROM3[7468]<=26'd9739101; ROM4[7468]<=26'd23458488;
ROM1[7469]<=26'd1968792; ROM2[7469]<=26'd11129572; ROM3[7469]<=26'd9747141; ROM4[7469]<=26'd23464829;
ROM1[7470]<=26'd1972791; ROM2[7470]<=26'd11138000; ROM3[7470]<=26'd9757002; ROM4[7470]<=26'd23474109;
ROM1[7471]<=26'd1964438; ROM2[7471]<=26'd11130716; ROM3[7471]<=26'd9747951; ROM4[7471]<=26'd23464621;
ROM1[7472]<=26'd1967163; ROM2[7472]<=26'd11125602; ROM3[7472]<=26'd9737789; ROM4[7472]<=26'd23457169;
ROM1[7473]<=26'd1975008; ROM2[7473]<=26'd11122261; ROM3[7473]<=26'd9729257; ROM4[7473]<=26'd23453760;
ROM1[7474]<=26'd1972787; ROM2[7474]<=26'd11119837; ROM3[7474]<=26'd9725370; ROM4[7474]<=26'd23452168;
ROM1[7475]<=26'd1975452; ROM2[7475]<=26'd11127992; ROM3[7475]<=26'd9733515; ROM4[7475]<=26'd23458197;
ROM1[7476]<=26'd1970785; ROM2[7476]<=26'd11130183; ROM3[7476]<=26'd9738474; ROM4[7476]<=26'd23461997;
ROM1[7477]<=26'd1961142; ROM2[7477]<=26'd11126392; ROM3[7477]<=26'd9737185; ROM4[7477]<=26'd23459706;
ROM1[7478]<=26'd1953581; ROM2[7478]<=26'd11124593; ROM3[7478]<=26'd9734608; ROM4[7478]<=26'd23456331;
ROM1[7479]<=26'd1952218; ROM2[7479]<=26'd11123864; ROM3[7479]<=26'd9733204; ROM4[7479]<=26'd23455707;
ROM1[7480]<=26'd1959722; ROM2[7480]<=26'd11125382; ROM3[7480]<=26'd9731964; ROM4[7480]<=26'd23454536;
ROM1[7481]<=26'd1972188; ROM2[7481]<=26'd11127508; ROM3[7481]<=26'd9725919; ROM4[7481]<=26'd23452224;
ROM1[7482]<=26'd1977294; ROM2[7482]<=26'd11124590; ROM3[7482]<=26'd9720821; ROM4[7482]<=26'd23449822;
ROM1[7483]<=26'd1974306; ROM2[7483]<=26'd11125543; ROM3[7483]<=26'd9722877; ROM4[7483]<=26'd23453374;
ROM1[7484]<=26'd1969502; ROM2[7484]<=26'd11129663; ROM3[7484]<=26'd9728636; ROM4[7484]<=26'd23457436;
ROM1[7485]<=26'd1967019; ROM2[7485]<=26'd11133947; ROM3[7485]<=26'd9735180; ROM4[7485]<=26'd23461490;
ROM1[7486]<=26'd1961616; ROM2[7486]<=26'd11134290; ROM3[7486]<=26'd9736098; ROM4[7486]<=26'd23460920;
ROM1[7487]<=26'd1962416; ROM2[7487]<=26'd11136438; ROM3[7487]<=26'd9740059; ROM4[7487]<=26'd23462032;
ROM1[7488]<=26'd1969417; ROM2[7488]<=26'd11138422; ROM3[7488]<=26'd9740932; ROM4[7488]<=26'd23463160;
ROM1[7489]<=26'd1972681; ROM2[7489]<=26'd11130272; ROM3[7489]<=26'd9728838; ROM4[7489]<=26'd23453533;
ROM1[7490]<=26'd1977439; ROM2[7490]<=26'd11124460; ROM3[7490]<=26'd9721424; ROM4[7490]<=26'd23448757;
ROM1[7491]<=26'd1973343; ROM2[7491]<=26'd11124408; ROM3[7491]<=26'd9720689; ROM4[7491]<=26'd23449475;
ROM1[7492]<=26'd1970214; ROM2[7492]<=26'd11127503; ROM3[7492]<=26'd9726087; ROM4[7492]<=26'd23453775;
ROM1[7493]<=26'd1972517; ROM2[7493]<=26'd11133436; ROM3[7493]<=26'd9736216; ROM4[7493]<=26'd23461995;
ROM1[7494]<=26'd1969291; ROM2[7494]<=26'd11135700; ROM3[7494]<=26'd9739950; ROM4[7494]<=26'd23462605;
ROM1[7495]<=26'd1960746; ROM2[7495]<=26'd11130659; ROM3[7495]<=26'd9738092; ROM4[7495]<=26'd23457334;
ROM1[7496]<=26'd1954768; ROM2[7496]<=26'd11124738; ROM3[7496]<=26'd9731454; ROM4[7496]<=26'd23451304;
ROM1[7497]<=26'd1958165; ROM2[7497]<=26'd11121571; ROM3[7497]<=26'd9724101; ROM4[7497]<=26'd23445960;
ROM1[7498]<=26'd1970098; ROM2[7498]<=26'd11121322; ROM3[7498]<=26'd9717560; ROM4[7498]<=26'd23444091;
ROM1[7499]<=26'd1974139; ROM2[7499]<=26'd11122192; ROM3[7499]<=26'd9717024; ROM4[7499]<=26'd23444845;
ROM1[7500]<=26'd1974773; ROM2[7500]<=26'd11128043; ROM3[7500]<=26'd9723684; ROM4[7500]<=26'd23450160;
ROM1[7501]<=26'd1972750; ROM2[7501]<=26'd11133324; ROM3[7501]<=26'd9731222; ROM4[7501]<=26'd23454755;
ROM1[7502]<=26'd1965182; ROM2[7502]<=26'd11132335; ROM3[7502]<=26'd9733330; ROM4[7502]<=26'd23454158;
ROM1[7503]<=26'd1958034; ROM2[7503]<=26'd11129873; ROM3[7503]<=26'd9735501; ROM4[7503]<=26'd23453496;
ROM1[7504]<=26'd1953418; ROM2[7504]<=26'd11125841; ROM3[7504]<=26'd9734870; ROM4[7504]<=26'd23452381;
ROM1[7505]<=26'd1959943; ROM2[7505]<=26'd11124202; ROM3[7505]<=26'd9732401; ROM4[7505]<=26'd23452435;
ROM1[7506]<=26'd1975100; ROM2[7506]<=26'd11126386; ROM3[7506]<=26'd9729428; ROM4[7506]<=26'd23454790;
ROM1[7507]<=26'd1986398; ROM2[7507]<=26'd11133228; ROM3[7507]<=26'd9731876; ROM4[7507]<=26'd23462662;
ROM1[7508]<=26'd1982649; ROM2[7508]<=26'd11134037; ROM3[7508]<=26'd9733525; ROM4[7508]<=26'd23463350;
ROM1[7509]<=26'd1967525; ROM2[7509]<=26'd11126075; ROM3[7509]<=26'd9731185; ROM4[7509]<=26'd23455995;
ROM1[7510]<=26'd1962968; ROM2[7510]<=26'd11126527; ROM3[7510]<=26'd9735719; ROM4[7510]<=26'd23458833;
ROM1[7511]<=26'd1958385; ROM2[7511]<=26'd11126178; ROM3[7511]<=26'd9738372; ROM4[7511]<=26'd23460661;
ROM1[7512]<=26'd1952526; ROM2[7512]<=26'd11124103; ROM3[7512]<=26'd9737245; ROM4[7512]<=26'd23458012;
ROM1[7513]<=26'd1956736; ROM2[7513]<=26'd11125845; ROM3[7513]<=26'd9735488; ROM4[7513]<=26'd23458458;
ROM1[7514]<=26'd1972190; ROM2[7514]<=26'd11133039; ROM3[7514]<=26'd9735332; ROM4[7514]<=26'd23462376;
ROM1[7515]<=26'd1982353; ROM2[7515]<=26'd11135015; ROM3[7515]<=26'd9730488; ROM4[7515]<=26'd23459939;
ROM1[7516]<=26'd1978721; ROM2[7516]<=26'd11132488; ROM3[7516]<=26'd9727602; ROM4[7516]<=26'd23456701;
ROM1[7517]<=26'd1973936; ROM2[7517]<=26'd11134027; ROM3[7517]<=26'd9732347; ROM4[7517]<=26'd23458261;
ROM1[7518]<=26'd1965341; ROM2[7518]<=26'd11128730; ROM3[7518]<=26'd9731784; ROM4[7518]<=26'd23453975;
ROM1[7519]<=26'd1963863; ROM2[7519]<=26'd11130564; ROM3[7519]<=26'd9737096; ROM4[7519]<=26'd23458586;
ROM1[7520]<=26'd1960823; ROM2[7520]<=26'd11132526; ROM3[7520]<=26'd9740721; ROM4[7520]<=26'd23460377;
ROM1[7521]<=26'd1954010; ROM2[7521]<=26'd11124320; ROM3[7521]<=26'd9731965; ROM4[7521]<=26'd23451677;
ROM1[7522]<=26'd1960847; ROM2[7522]<=26'd11124002; ROM3[7522]<=26'd9727580; ROM4[7522]<=26'd23450164;
ROM1[7523]<=26'd1971202; ROM2[7523]<=26'd11122914; ROM3[7523]<=26'd9720208; ROM4[7523]<=26'd23447555;
ROM1[7524]<=26'd1975903; ROM2[7524]<=26'd11123252; ROM3[7524]<=26'd9720310; ROM4[7524]<=26'd23449407;
ROM1[7525]<=26'd1979785; ROM2[7525]<=26'd11132799; ROM3[7525]<=26'd9731678; ROM4[7525]<=26'd23460941;
ROM1[7526]<=26'd1973358; ROM2[7526]<=26'd11133489; ROM3[7526]<=26'd9735850; ROM4[7526]<=26'd23463117;
ROM1[7527]<=26'd1962782; ROM2[7527]<=26'd11127135; ROM3[7527]<=26'd9733758; ROM4[7527]<=26'd23457387;
ROM1[7528]<=26'd1955616; ROM2[7528]<=26'd11125127; ROM3[7528]<=26'd9735288; ROM4[7528]<=26'd23457114;
ROM1[7529]<=26'd1956294; ROM2[7529]<=26'd11126505; ROM3[7529]<=26'd9738510; ROM4[7529]<=26'd23459046;
ROM1[7530]<=26'd1964017; ROM2[7530]<=26'd11128867; ROM3[7530]<=26'd9738598; ROM4[7530]<=26'd23460485;
ROM1[7531]<=26'd1974314; ROM2[7531]<=26'd11128657; ROM3[7531]<=26'd9732106; ROM4[7531]<=26'd23459271;
ROM1[7532]<=26'd1981039; ROM2[7532]<=26'd11127878; ROM3[7532]<=26'd9728831; ROM4[7532]<=26'd23457738;
ROM1[7533]<=26'd1979834; ROM2[7533]<=26'd11130157; ROM3[7533]<=26'd9733090; ROM4[7533]<=26'd23460231;
ROM1[7534]<=26'd1974624; ROM2[7534]<=26'd11132079; ROM3[7534]<=26'd9736883; ROM4[7534]<=26'd23462533;
ROM1[7535]<=26'd1968243; ROM2[7535]<=26'd11130100; ROM3[7535]<=26'd9737871; ROM4[7535]<=26'd23461378;
ROM1[7536]<=26'd1966043; ROM2[7536]<=26'd11132970; ROM3[7536]<=26'd9743458; ROM4[7536]<=26'd23465610;
ROM1[7537]<=26'd1973132; ROM2[7537]<=26'd11141565; ROM3[7537]<=26'd9752873; ROM4[7537]<=26'd23473536;
ROM1[7538]<=26'd1974870; ROM2[7538]<=26'd11137001; ROM3[7538]<=26'd9748653; ROM4[7538]<=26'd23468959;
ROM1[7539]<=26'd1979528; ROM2[7539]<=26'd11132074; ROM3[7539]<=26'd9740034; ROM4[7539]<=26'd23463051;
ROM1[7540]<=26'd1985378; ROM2[7540]<=26'd11128861; ROM3[7540]<=26'd9730039; ROM4[7540]<=26'd23457618;
ROM1[7541]<=26'd1979648; ROM2[7541]<=26'd11124202; ROM3[7541]<=26'd9724806; ROM4[7541]<=26'd23452326;
ROM1[7542]<=26'd1979248; ROM2[7542]<=26'd11131316; ROM3[7542]<=26'd9733692; ROM4[7542]<=26'd23458687;
ROM1[7543]<=26'd1977943; ROM2[7543]<=26'd11135200; ROM3[7543]<=26'd9740206; ROM4[7543]<=26'd23463068;
ROM1[7544]<=26'd1967689; ROM2[7544]<=26'd11128517; ROM3[7544]<=26'd9738915; ROM4[7544]<=26'd23457767;
ROM1[7545]<=26'd1955444; ROM2[7545]<=26'd11121951; ROM3[7545]<=26'd9735383; ROM4[7545]<=26'd23451667;
ROM1[7546]<=26'd1953251; ROM2[7546]<=26'd11120968; ROM3[7546]<=26'd9730358; ROM4[7546]<=26'd23448344;
ROM1[7547]<=26'd1964789; ROM2[7547]<=26'd11127634; ROM3[7547]<=26'd9730190; ROM4[7547]<=26'd23452850;
ROM1[7548]<=26'd1980924; ROM2[7548]<=26'd11134164; ROM3[7548]<=26'd9729979; ROM4[7548]<=26'd23456363;
ROM1[7549]<=26'd1981796; ROM2[7549]<=26'd11131305; ROM3[7549]<=26'd9726578; ROM4[7549]<=26'd23452939;
ROM1[7550]<=26'd1974872; ROM2[7550]<=26'd11126093; ROM3[7550]<=26'd9726622; ROM4[7550]<=26'd23449313;
ROM1[7551]<=26'd1967212; ROM2[7551]<=26'd11124051; ROM3[7551]<=26'd9729065; ROM4[7551]<=26'd23447541;
ROM1[7552]<=26'd1963007; ROM2[7552]<=26'd11125255; ROM3[7552]<=26'd9732096; ROM4[7552]<=26'd23449481;
ROM1[7553]<=26'd1957862; ROM2[7553]<=26'd11124610; ROM3[7553]<=26'd9733861; ROM4[7553]<=26'd23451525;
ROM1[7554]<=26'd1956485; ROM2[7554]<=26'd11124126; ROM3[7554]<=26'd9735410; ROM4[7554]<=26'd23453226;
ROM1[7555]<=26'd1965335; ROM2[7555]<=26'd11125690; ROM3[7555]<=26'd9734628; ROM4[7555]<=26'd23453059;
ROM1[7556]<=26'd1982187; ROM2[7556]<=26'd11129789; ROM3[7556]<=26'd9732386; ROM4[7556]<=26'd23455538;
ROM1[7557]<=26'd1993022; ROM2[7557]<=26'd11135292; ROM3[7557]<=26'd9733628; ROM4[7557]<=26'd23460536;
ROM1[7558]<=26'd1989158; ROM2[7558]<=26'd11135104; ROM3[7558]<=26'd9733895; ROM4[7558]<=26'd23461184;
ROM1[7559]<=26'd1982569; ROM2[7559]<=26'd11132742; ROM3[7559]<=26'd9736464; ROM4[7559]<=26'd23459798;
ROM1[7560]<=26'd1979364; ROM2[7560]<=26'd11135521; ROM3[7560]<=26'd9742626; ROM4[7560]<=26'd23464717;
ROM1[7561]<=26'd1977340; ROM2[7561]<=26'd11140012; ROM3[7561]<=26'd9750743; ROM4[7561]<=26'd23469548;
ROM1[7562]<=26'd1964972; ROM2[7562]<=26'd11131052; ROM3[7562]<=26'd9743137; ROM4[7562]<=26'd23458475;
ROM1[7563]<=26'd1958776; ROM2[7563]<=26'd11122820; ROM3[7563]<=26'd9730133; ROM4[7563]<=26'd23448603;
ROM1[7564]<=26'd1966246; ROM2[7564]<=26'd11118865; ROM3[7564]<=26'd9722143; ROM4[7564]<=26'd23442539;
ROM1[7565]<=26'd1970853; ROM2[7565]<=26'd11113941; ROM3[7565]<=26'd9711342; ROM4[7565]<=26'd23436931;
ROM1[7566]<=26'd1972545; ROM2[7566]<=26'd11119138; ROM3[7566]<=26'd9715596; ROM4[7566]<=26'd23442933;
ROM1[7567]<=26'd1970480; ROM2[7567]<=26'd11123342; ROM3[7567]<=26'd9724402; ROM4[7567]<=26'd23448902;
ROM1[7568]<=26'd1963287; ROM2[7568]<=26'd11122790; ROM3[7568]<=26'd9727760; ROM4[7568]<=26'd23450115;
ROM1[7569]<=26'd1956384; ROM2[7569]<=26'd11121538; ROM3[7569]<=26'd9727977; ROM4[7569]<=26'd23448443;
ROM1[7570]<=26'd1953590; ROM2[7570]<=26'd11122680; ROM3[7570]<=26'd9730209; ROM4[7570]<=26'd23450075;
ROM1[7571]<=26'd1957807; ROM2[7571]<=26'd11124874; ROM3[7571]<=26'd9732620; ROM4[7571]<=26'd23453300;
ROM1[7572]<=26'd1966330; ROM2[7572]<=26'd11126826; ROM3[7572]<=26'd9729520; ROM4[7572]<=26'd23453139;
ROM1[7573]<=26'd1984672; ROM2[7573]<=26'd11134707; ROM3[7573]<=26'd9730083; ROM4[7573]<=26'd23458261;
ROM1[7574]<=26'd1993377; ROM2[7574]<=26'd11140529; ROM3[7574]<=26'd9734888; ROM4[7574]<=26'd23462357;
ROM1[7575]<=26'd1984574; ROM2[7575]<=26'd11138668; ROM3[7575]<=26'd9733798; ROM4[7575]<=26'd23459480;
ROM1[7576]<=26'd1970303; ROM2[7576]<=26'd11131956; ROM3[7576]<=26'd9729524; ROM4[7576]<=26'd23455302;
ROM1[7577]<=26'd1958351; ROM2[7577]<=26'd11124216; ROM3[7577]<=26'd9727292; ROM4[7577]<=26'd23450134;
ROM1[7578]<=26'd1951319; ROM2[7578]<=26'd11121059; ROM3[7578]<=26'd9729866; ROM4[7578]<=26'd23449398;
ROM1[7579]<=26'd1953518; ROM2[7579]<=26'd11122778; ROM3[7579]<=26'd9733893; ROM4[7579]<=26'd23452555;
ROM1[7580]<=26'd1964355; ROM2[7580]<=26'd11125880; ROM3[7580]<=26'd9734154; ROM4[7580]<=26'd23453789;
ROM1[7581]<=26'd1979631; ROM2[7581]<=26'd11129896; ROM3[7581]<=26'd9732311; ROM4[7581]<=26'd23456461;
ROM1[7582]<=26'd1986305; ROM2[7582]<=26'd11130791; ROM3[7582]<=26'd9730657; ROM4[7582]<=26'd23458423;
ROM1[7583]<=26'd1984321; ROM2[7583]<=26'd11132337; ROM3[7583]<=26'd9735044; ROM4[7583]<=26'd23460169;
ROM1[7584]<=26'd1981507; ROM2[7584]<=26'd11136180; ROM3[7584]<=26'd9742755; ROM4[7584]<=26'd23463711;
ROM1[7585]<=26'd1975583; ROM2[7585]<=26'd11134186; ROM3[7585]<=26'd9743278; ROM4[7585]<=26'd23462637;
ROM1[7586]<=26'd1969987; ROM2[7586]<=26'd11133814; ROM3[7586]<=26'd9745021; ROM4[7586]<=26'd23461841;
ROM1[7587]<=26'd1973361; ROM2[7587]<=26'd11140902; ROM3[7587]<=26'd9752324; ROM4[7587]<=26'd23468224;
ROM1[7588]<=26'd1980398; ROM2[7588]<=26'd11145273; ROM3[7588]<=26'd9752700; ROM4[7588]<=26'd23470713;
ROM1[7589]<=26'd1990331; ROM2[7589]<=26'd11145372; ROM3[7589]<=26'd9746188; ROM4[7589]<=26'd23467300;
ROM1[7590]<=26'd2002820; ROM2[7590]<=26'd11147688; ROM3[7590]<=26'd9743223; ROM4[7590]<=26'd23469350;
ROM1[7591]<=26'd2002684; ROM2[7591]<=26'd11148377; ROM3[7591]<=26'd9743648; ROM4[7591]<=26'd23469464;
ROM1[7592]<=26'd1995164; ROM2[7592]<=26'd11144088; ROM3[7592]<=26'd9742891; ROM4[7592]<=26'd23467181;
ROM1[7593]<=26'd1988771; ROM2[7593]<=26'd11142993; ROM3[7593]<=26'd9746949; ROM4[7593]<=26'd23469382;
ROM1[7594]<=26'd1981105; ROM2[7594]<=26'd11142821; ROM3[7594]<=26'd9748407; ROM4[7594]<=26'd23468285;
ROM1[7595]<=26'd1971645; ROM2[7595]<=26'd11137524; ROM3[7595]<=26'd9746780; ROM4[7595]<=26'd23464378;
ROM1[7596]<=26'd1971206; ROM2[7596]<=26'd11134642; ROM3[7596]<=26'd9745917; ROM4[7596]<=26'd23463909;
ROM1[7597]<=26'd1982196; ROM2[7597]<=26'd11137052; ROM3[7597]<=26'd9742091; ROM4[7597]<=26'd23463845;
ROM1[7598]<=26'd1994935; ROM2[7598]<=26'd11138962; ROM3[7598]<=26'd9736820; ROM4[7598]<=26'd23462309;
ROM1[7599]<=26'd1998377; ROM2[7599]<=26'd11139995; ROM3[7599]<=26'd9735940; ROM4[7599]<=26'd23464357;
ROM1[7600]<=26'd1996502; ROM2[7600]<=26'd11145438; ROM3[7600]<=26'd9743536; ROM4[7600]<=26'd23469099;
ROM1[7601]<=26'd1993409; ROM2[7601]<=26'd11149500; ROM3[7601]<=26'd9750662; ROM4[7601]<=26'd23471663;
ROM1[7602]<=26'd1989376; ROM2[7602]<=26'd11147690; ROM3[7602]<=26'd9752507; ROM4[7602]<=26'd23472586;
ROM1[7603]<=26'd1979254; ROM2[7603]<=26'd11141875; ROM3[7603]<=26'd9749862; ROM4[7603]<=26'd23467362;
ROM1[7604]<=26'd1982809; ROM2[7604]<=26'd11146254; ROM3[7604]<=26'd9752920; ROM4[7604]<=26'd23469217;
ROM1[7605]<=26'd1994768; ROM2[7605]<=26'd11152441; ROM3[7605]<=26'd9755261; ROM4[7605]<=26'd23474915;
ROM1[7606]<=26'd1999538; ROM2[7606]<=26'd11144565; ROM3[7606]<=26'd9741758; ROM4[7606]<=26'd23464866;
ROM1[7607]<=26'd1998764; ROM2[7607]<=26'd11139136; ROM3[7607]<=26'd9732327; ROM4[7607]<=26'd23457272;
ROM1[7608]<=26'd1989981; ROM2[7608]<=26'd11134684; ROM3[7608]<=26'd9730517; ROM4[7608]<=26'd23455402;
ROM1[7609]<=26'd1975638; ROM2[7609]<=26'd11128083; ROM3[7609]<=26'd9726611; ROM4[7609]<=26'd23447466;
ROM1[7610]<=26'd1970795; ROM2[7610]<=26'd11129914; ROM3[7610]<=26'd9728871; ROM4[7610]<=26'd23448759;
ROM1[7611]<=26'd1970164; ROM2[7611]<=26'd11134420; ROM3[7611]<=26'd9735436; ROM4[7611]<=26'd23454765;
ROM1[7612]<=26'd1966676; ROM2[7612]<=26'd11134092; ROM3[7612]<=26'd9734212; ROM4[7612]<=26'd23453147;
ROM1[7613]<=26'd1968146; ROM2[7613]<=26'd11131250; ROM3[7613]<=26'd9729844; ROM4[7613]<=26'd23450699;
ROM1[7614]<=26'd1978825; ROM2[7614]<=26'd11130851; ROM3[7614]<=26'd9727023; ROM4[7614]<=26'd23449891;
ROM1[7615]<=26'd1988791; ROM2[7615]<=26'd11132332; ROM3[7615]<=26'd9722991; ROM4[7615]<=26'd23449227;
ROM1[7616]<=26'd1987114; ROM2[7616]<=26'd11133802; ROM3[7616]<=26'd9723906; ROM4[7616]<=26'd23450776;
ROM1[7617]<=26'd1978430; ROM2[7617]<=26'd11132494; ROM3[7617]<=26'd9725594; ROM4[7617]<=26'd23451094;
ROM1[7618]<=26'd1974430; ROM2[7618]<=26'd11135169; ROM3[7618]<=26'd9732717; ROM4[7618]<=26'd23455411;
ROM1[7619]<=26'd1976973; ROM2[7619]<=26'd11141831; ROM3[7619]<=26'd9744586; ROM4[7619]<=26'd23465230;
ROM1[7620]<=26'd1969056; ROM2[7620]<=26'd11136510; ROM3[7620]<=26'd9745493; ROM4[7620]<=26'd23462381;
ROM1[7621]<=26'd1964852; ROM2[7621]<=26'd11129932; ROM3[7621]<=26'd9741175; ROM4[7621]<=26'd23456733;
ROM1[7622]<=26'd1973619; ROM2[7622]<=26'd11130378; ROM3[7622]<=26'd9739474; ROM4[7622]<=26'd23457106;
ROM1[7623]<=26'd1985252; ROM2[7623]<=26'd11132523; ROM3[7623]<=26'd9734282; ROM4[7623]<=26'd23457163;
ROM1[7624]<=26'd1985411; ROM2[7624]<=26'd11130588; ROM3[7624]<=26'd9731105; ROM4[7624]<=26'd23454369;
ROM1[7625]<=26'd1982345; ROM2[7625]<=26'd11131388; ROM3[7625]<=26'd9737360; ROM4[7625]<=26'd23457621;
ROM1[7626]<=26'd1982286; ROM2[7626]<=26'd11137559; ROM3[7626]<=26'd9744652; ROM4[7626]<=26'd23463798;
ROM1[7627]<=26'd1979974; ROM2[7627]<=26'd11139864; ROM3[7627]<=26'd9746529; ROM4[7627]<=26'd23464744;
ROM1[7628]<=26'd1965867; ROM2[7628]<=26'd11132940; ROM3[7628]<=26'd9740770; ROM4[7628]<=26'd23458045;
ROM1[7629]<=26'd1959594; ROM2[7629]<=26'd11129790; ROM3[7629]<=26'd9735422; ROM4[7629]<=26'd23454379;
ROM1[7630]<=26'd1968006; ROM2[7630]<=26'd11131576; ROM3[7630]<=26'd9732577; ROM4[7630]<=26'd23456001;
ROM1[7631]<=26'd1983457; ROM2[7631]<=26'd11133404; ROM3[7631]<=26'd9729822; ROM4[7631]<=26'd23458637;
ROM1[7632]<=26'd1999709; ROM2[7632]<=26'd11141677; ROM3[7632]<=26'd9733942; ROM4[7632]<=26'd23466313;
ROM1[7633]<=26'd2001729; ROM2[7633]<=26'd11146636; ROM3[7633]<=26'd9738578; ROM4[7633]<=26'd23471134;
ROM1[7634]<=26'd1988406; ROM2[7634]<=26'd11143741; ROM3[7634]<=26'd9738940; ROM4[7634]<=26'd23468845;
ROM1[7635]<=26'd1979749; ROM2[7635]<=26'd11139418; ROM3[7635]<=26'd9739502; ROM4[7635]<=26'd23464947;
ROM1[7636]<=26'd1977926; ROM2[7636]<=26'd11140184; ROM3[7636]<=26'd9741391; ROM4[7636]<=26'd23466421;
ROM1[7637]<=26'd1976509; ROM2[7637]<=26'd11143967; ROM3[7637]<=26'd9743696; ROM4[7637]<=26'd23468784;
ROM1[7638]<=26'd1985813; ROM2[7638]<=26'd11146962; ROM3[7638]<=26'd9742524; ROM4[7638]<=26'd23469299;
ROM1[7639]<=26'd2005894; ROM2[7639]<=26'd11153705; ROM3[7639]<=26'd9742592; ROM4[7639]<=26'd23475130;
ROM1[7640]<=26'd2018475; ROM2[7640]<=26'd11157928; ROM3[7640]<=26'd9745502; ROM4[7640]<=26'd23480019;
ROM1[7641]<=26'd2013326; ROM2[7641]<=26'd11157384; ROM3[7641]<=26'd9747743; ROM4[7641]<=26'd23479429;
ROM1[7642]<=26'd2007143; ROM2[7642]<=26'd11157678; ROM3[7642]<=26'd9751416; ROM4[7642]<=26'd23480995;
ROM1[7643]<=26'd1995892; ROM2[7643]<=26'd11151239; ROM3[7643]<=26'd9747749; ROM4[7643]<=26'd23474874;
ROM1[7644]<=26'd1993196; ROM2[7644]<=26'd11153354; ROM3[7644]<=26'd9747323; ROM4[7644]<=26'd23473271;
ROM1[7645]<=26'd1990677; ROM2[7645]<=26'd11153369; ROM3[7645]<=26'd9750816; ROM4[7645]<=26'd23473432;
ROM1[7646]<=26'd1989504; ROM2[7646]<=26'd11152370; ROM3[7646]<=26'd9752330; ROM4[7646]<=26'd23473043;
ROM1[7647]<=26'd2019223; ROM2[7647]<=26'd11166680; ROM3[7647]<=26'd9759780; ROM4[7647]<=26'd23485347;
ROM1[7648]<=26'd2036031; ROM2[7648]<=26'd11168526; ROM3[7648]<=26'd9756325; ROM4[7648]<=26'd23487023;
ROM1[7649]<=26'd2043266; ROM2[7649]<=26'd11170218; ROM3[7649]<=26'd9752547; ROM4[7649]<=26'd23486865;
ROM1[7650]<=26'd2045667; ROM2[7650]<=26'd11168983; ROM3[7650]<=26'd9756316; ROM4[7650]<=26'd23489031;
ROM1[7651]<=26'd2032545; ROM2[7651]<=26'd11161567; ROM3[7651]<=26'd9756824; ROM4[7651]<=26'd23484482;
ROM1[7652]<=26'd2036142; ROM2[7652]<=26'd11164400; ROM3[7652]<=26'd9762551; ROM4[7652]<=26'd23488861;
ROM1[7653]<=26'd2044817; ROM2[7653]<=26'd11168853; ROM3[7653]<=26'd9770900; ROM4[7653]<=26'd23496034;
ROM1[7654]<=26'd2055887; ROM2[7654]<=26'd11175281; ROM3[7654]<=26'd9771408; ROM4[7654]<=26'd23498102;
ROM1[7655]<=26'd2069552; ROM2[7655]<=26'd11180841; ROM3[7655]<=26'd9769050; ROM4[7655]<=26'd23500182;
ROM1[7656]<=26'd2091575; ROM2[7656]<=26'd11186630; ROM3[7656]<=26'd9768816; ROM4[7656]<=26'd23504213;
ROM1[7657]<=26'd2108860; ROM2[7657]<=26'd11192059; ROM3[7657]<=26'd9769951; ROM4[7657]<=26'd23509208;
ROM1[7658]<=26'd2118505; ROM2[7658]<=26'd11198795; ROM3[7658]<=26'd9776623; ROM4[7658]<=26'd23515356;
ROM1[7659]<=26'd2116603; ROM2[7659]<=26'd11198262; ROM3[7659]<=26'd9778122; ROM4[7659]<=26'd23514003;
ROM1[7660]<=26'd2119670; ROM2[7660]<=26'd11201325; ROM3[7660]<=26'd9780487; ROM4[7660]<=26'd23514169;
ROM1[7661]<=26'd2135918; ROM2[7661]<=26'd11211641; ROM3[7661]<=26'd9792039; ROM4[7661]<=26'd23523501;
ROM1[7662]<=26'd2138988; ROM2[7662]<=26'd11210171; ROM3[7662]<=26'd9791233; ROM4[7662]<=26'd23523224;
ROM1[7663]<=26'd2139979; ROM2[7663]<=26'd11204317; ROM3[7663]<=26'd9782637; ROM4[7663]<=26'd23515017;
ROM1[7664]<=26'd2153432; ROM2[7664]<=26'd11201426; ROM3[7664]<=26'd9774653; ROM4[7664]<=26'd23510019;
ROM1[7665]<=26'd2165955; ROM2[7665]<=26'd11200351; ROM3[7665]<=26'd9767648; ROM4[7665]<=26'd23508698;
ROM1[7666]<=26'd2170743; ROM2[7666]<=26'd11202822; ROM3[7666]<=26'd9767327; ROM4[7666]<=26'd23509795;
ROM1[7667]<=26'd2178689; ROM2[7667]<=26'd11210390; ROM3[7667]<=26'd9774005; ROM4[7667]<=26'd23516587;
ROM1[7668]<=26'd2179477; ROM2[7668]<=26'd11212540; ROM3[7668]<=26'd9777593; ROM4[7668]<=26'd23520267;
ROM1[7669]<=26'd2173645; ROM2[7669]<=26'd11210226; ROM3[7669]<=26'd9775770; ROM4[7669]<=26'd23518157;
ROM1[7670]<=26'd2170599; ROM2[7670]<=26'd11210029; ROM3[7670]<=26'd9778188; ROM4[7670]<=26'd23517536;
ROM1[7671]<=26'd2176620; ROM2[7671]<=26'd11213520; ROM3[7671]<=26'd9780048; ROM4[7671]<=26'd23519168;
ROM1[7672]<=26'd2191313; ROM2[7672]<=26'd11216962; ROM3[7672]<=26'd9776677; ROM4[7672]<=26'd23520395;
ROM1[7673]<=26'd2210994; ROM2[7673]<=26'd11222276; ROM3[7673]<=26'd9773725; ROM4[7673]<=26'd23523647;
ROM1[7674]<=26'd2225773; ROM2[7674]<=26'd11233364; ROM3[7674]<=26'd9782388; ROM4[7674]<=26'd23535203;
ROM1[7675]<=26'd2234145; ROM2[7675]<=26'd11242353; ROM3[7675]<=26'd9793511; ROM4[7675]<=26'd23546728;
ROM1[7676]<=26'd2227776; ROM2[7676]<=26'd11239805; ROM3[7676]<=26'd9794408; ROM4[7676]<=26'd23546294;
ROM1[7677]<=26'd2226613; ROM2[7677]<=26'd11243223; ROM3[7677]<=26'd9798826; ROM4[7677]<=26'd23548686;
ROM1[7678]<=26'd2226482; ROM2[7678]<=26'd11245379; ROM3[7678]<=26'd9801943; ROM4[7678]<=26'd23552011;
ROM1[7679]<=26'd2218982; ROM2[7679]<=26'd11233908; ROM3[7679]<=26'd9792176; ROM4[7679]<=26'd23544098;
ROM1[7680]<=26'd2227604; ROM2[7680]<=26'd11233419; ROM3[7680]<=26'd9790014; ROM4[7680]<=26'd23544187;
ROM1[7681]<=26'd2240132; ROM2[7681]<=26'd11234196; ROM3[7681]<=26'd9785771; ROM4[7681]<=26'd23545176;
ROM1[7682]<=26'd2244782; ROM2[7682]<=26'd11231806; ROM3[7682]<=26'd9781094; ROM4[7682]<=26'd23542088;
ROM1[7683]<=26'd2244653; ROM2[7683]<=26'd11236001; ROM3[7683]<=26'd9788664; ROM4[7683]<=26'd23546311;
ROM1[7684]<=26'd2247281; ROM2[7684]<=26'd11244570; ROM3[7684]<=26'd9799361; ROM4[7684]<=26'd23553491;
ROM1[7685]<=26'd2242513; ROM2[7685]<=26'd11242366; ROM3[7685]<=26'd9801119; ROM4[7685]<=26'd23552393;
ROM1[7686]<=26'd2229422; ROM2[7686]<=26'd11233714; ROM3[7686]<=26'd9794709; ROM4[7686]<=26'd23545368;
ROM1[7687]<=26'd2224459; ROM2[7687]<=26'd11231979; ROM3[7687]<=26'd9795046; ROM4[7687]<=26'd23542907;
ROM1[7688]<=26'd2228421; ROM2[7688]<=26'd11232919; ROM3[7688]<=26'd9797264; ROM4[7688]<=26'd23545779;
ROM1[7689]<=26'd2238115; ROM2[7689]<=26'd11231448; ROM3[7689]<=26'd9791749; ROM4[7689]<=26'd23544746;
ROM1[7690]<=26'd2250203; ROM2[7690]<=26'd11233287; ROM3[7690]<=26'd9790265; ROM4[7690]<=26'd23546160;
ROM1[7691]<=26'd2249110; ROM2[7691]<=26'd11233704; ROM3[7691]<=26'd9792756; ROM4[7691]<=26'd23549697;
ROM1[7692]<=26'd2237233; ROM2[7692]<=26'd11230571; ROM3[7692]<=26'd9792845; ROM4[7692]<=26'd23547019;
ROM1[7693]<=26'd2228980; ROM2[7693]<=26'd11229616; ROM3[7693]<=26'd9796098; ROM4[7693]<=26'd23546440;
ROM1[7694]<=26'd2221455; ROM2[7694]<=26'd11228222; ROM3[7694]<=26'd9796137; ROM4[7694]<=26'd23545848;
ROM1[7695]<=26'd2214157; ROM2[7695]<=26'd11226616; ROM3[7695]<=26'd9794685; ROM4[7695]<=26'd23544635;
ROM1[7696]<=26'd2210889; ROM2[7696]<=26'd11224085; ROM3[7696]<=26'd9791506; ROM4[7696]<=26'd23542037;
ROM1[7697]<=26'd2216692; ROM2[7697]<=26'd11224216; ROM3[7697]<=26'd9786887; ROM4[7697]<=26'd23540267;
ROM1[7698]<=26'd2226974; ROM2[7698]<=26'd11225698; ROM3[7698]<=26'd9783639; ROM4[7698]<=26'd23539673;
ROM1[7699]<=26'd2226084; ROM2[7699]<=26'd11228879; ROM3[7699]<=26'd9783959; ROM4[7699]<=26'd23541473;
ROM1[7700]<=26'd2223181; ROM2[7700]<=26'd11233847; ROM3[7700]<=26'd9790638; ROM4[7700]<=26'd23547751;
ROM1[7701]<=26'd2210602; ROM2[7701]<=26'd11228901; ROM3[7701]<=26'd9792641; ROM4[7701]<=26'd23544744;
ROM1[7702]<=26'd2195764; ROM2[7702]<=26'd11223071; ROM3[7702]<=26'd9792827; ROM4[7702]<=26'd23541399;
ROM1[7703]<=26'd2181046; ROM2[7703]<=26'd11216435; ROM3[7703]<=26'd9792492; ROM4[7703]<=26'd23536234;
ROM1[7704]<=26'd2168359; ROM2[7704]<=26'd11209309; ROM3[7704]<=26'd9787295; ROM4[7704]<=26'd23529213;
ROM1[7705]<=26'd2171699; ROM2[7705]<=26'd11210054; ROM3[7705]<=26'd9785256; ROM4[7705]<=26'd23530034;
ROM1[7706]<=26'd2181215; ROM2[7706]<=26'd11212954; ROM3[7706]<=26'd9783176; ROM4[7706]<=26'd23530870;
ROM1[7707]<=26'd2177611; ROM2[7707]<=26'd11207931; ROM3[7707]<=26'd9775637; ROM4[7707]<=26'd23526987;
ROM1[7708]<=26'd2163740; ROM2[7708]<=26'd11199304; ROM3[7708]<=26'd9772733; ROM4[7708]<=26'd23519976;
ROM1[7709]<=26'd2152438; ROM2[7709]<=26'd11196597; ROM3[7709]<=26'd9776642; ROM4[7709]<=26'd23519022;
ROM1[7710]<=26'd2142109; ROM2[7710]<=26'd11193975; ROM3[7710]<=26'd9775511; ROM4[7710]<=26'd23517721;
ROM1[7711]<=26'd2135924; ROM2[7711]<=26'd11195753; ROM3[7711]<=26'd9779986; ROM4[7711]<=26'd23517243;
ROM1[7712]<=26'd2137445; ROM2[7712]<=26'd11204300; ROM3[7712]<=26'd9787961; ROM4[7712]<=26'd23522826;
ROM1[7713]<=26'd2143429; ROM2[7713]<=26'd11211865; ROM3[7713]<=26'd9790258; ROM4[7713]<=26'd23526998;
ROM1[7714]<=26'd2149783; ROM2[7714]<=26'd11210336; ROM3[7714]<=26'd9785845; ROM4[7714]<=26'd23524330;
ROM1[7715]<=26'd2149112; ROM2[7715]<=26'd11200155; ROM3[7715]<=26'd9772025; ROM4[7715]<=26'd23514911;
ROM1[7716]<=26'd2136798; ROM2[7716]<=26'd11190875; ROM3[7716]<=26'd9764733; ROM4[7716]<=26'd23507395;
ROM1[7717]<=26'd2119852; ROM2[7717]<=26'd11183848; ROM3[7717]<=26'd9762043; ROM4[7717]<=26'd23501467;
ROM1[7718]<=26'd2108817; ROM2[7718]<=26'd11181128; ROM3[7718]<=26'd9764383; ROM4[7718]<=26'd23500960;
ROM1[7719]<=26'd2101925; ROM2[7719]<=26'd11180952; ROM3[7719]<=26'd9771024; ROM4[7719]<=26'd23502816;
ROM1[7720]<=26'd2089470; ROM2[7720]<=26'd11173517; ROM3[7720]<=26'd9769187; ROM4[7720]<=26'd23496579;
ROM1[7721]<=26'd2085152; ROM2[7721]<=26'd11169504; ROM3[7721]<=26'd9767757; ROM4[7721]<=26'd23493480;
ROM1[7722]<=26'd2093601; ROM2[7722]<=26'd11171434; ROM3[7722]<=26'd9765341; ROM4[7722]<=26'd23492728;
ROM1[7723]<=26'd2108739; ROM2[7723]<=26'd11177094; ROM3[7723]<=26'd9764136; ROM4[7723]<=26'd23495755;
ROM1[7724]<=26'd2108394; ROM2[7724]<=26'd11178017; ROM3[7724]<=26'd9763610; ROM4[7724]<=26'd23497979;
ROM1[7725]<=26'd2098883; ROM2[7725]<=26'd11175347; ROM3[7725]<=26'd9763570; ROM4[7725]<=26'd23496613;
ROM1[7726]<=26'd2092275; ROM2[7726]<=26'd11175254; ROM3[7726]<=26'd9769338; ROM4[7726]<=26'd23499474;
ROM1[7727]<=26'd2083563; ROM2[7727]<=26'd11172807; ROM3[7727]<=26'd9770995; ROM4[7727]<=26'd23498666;
ROM1[7728]<=26'd2070405; ROM2[7728]<=26'd11165721; ROM3[7728]<=26'd9765093; ROM4[7728]<=26'd23491523;
ROM1[7729]<=26'd2064153; ROM2[7729]<=26'd11161100; ROM3[7729]<=26'd9759297; ROM4[7729]<=26'd23485877;
ROM1[7730]<=26'd2066165; ROM2[7730]<=26'd11158793; ROM3[7730]<=26'd9752929; ROM4[7730]<=26'd23481765;
ROM1[7731]<=26'd2079288; ROM2[7731]<=26'd11162846; ROM3[7731]<=26'd9750448; ROM4[7731]<=26'd23485429;
ROM1[7732]<=26'd2093882; ROM2[7732]<=26'd11171939; ROM3[7732]<=26'd9757944; ROM4[7732]<=26'd23495121;
ROM1[7733]<=26'd2087047; ROM2[7733]<=26'd11167714; ROM3[7733]<=26'd9757857; ROM4[7733]<=26'd23492896;
ROM1[7734]<=26'd2073207; ROM2[7734]<=26'd11164395; ROM3[7734]<=26'd9757688; ROM4[7734]<=26'd23489892;
ROM1[7735]<=26'd2065556; ROM2[7735]<=26'd11165082; ROM3[7735]<=26'd9762228; ROM4[7735]<=26'd23493165;
ROM1[7736]<=26'd2058799; ROM2[7736]<=26'd11163455; ROM3[7736]<=26'd9765414; ROM4[7736]<=26'd23494680;
ROM1[7737]<=26'd2058527; ROM2[7737]<=26'd11167115; ROM3[7737]<=26'd9771906; ROM4[7737]<=26'd23498497;
ROM1[7738]<=26'd2063092; ROM2[7738]<=26'd11166655; ROM3[7738]<=26'd9771400; ROM4[7738]<=26'd23498641;
ROM1[7739]<=26'd2077991; ROM2[7739]<=26'd11170808; ROM3[7739]<=26'd9770248; ROM4[7739]<=26'd23501445;
ROM1[7740]<=26'd2091647; ROM2[7740]<=26'd11176397; ROM3[7740]<=26'd9772551; ROM4[7740]<=26'd23507798;
ROM1[7741]<=26'd2085274; ROM2[7741]<=26'd11173428; ROM3[7741]<=26'd9771302; ROM4[7741]<=26'd23507718;
ROM1[7742]<=26'd2071067; ROM2[7742]<=26'd11165569; ROM3[7742]<=26'd9768267; ROM4[7742]<=26'd23502586;
ROM1[7743]<=26'd2058838; ROM2[7743]<=26'd11158948; ROM3[7743]<=26'd9768224; ROM4[7743]<=26'd23496855;
ROM1[7744]<=26'd2047365; ROM2[7744]<=26'd11156388; ROM3[7744]<=26'd9766472; ROM4[7744]<=26'd23492853;
ROM1[7745]<=26'd2041328; ROM2[7745]<=26'd11155678; ROM3[7745]<=26'd9767500; ROM4[7745]<=26'd23492566;
ROM1[7746]<=26'd2047492; ROM2[7746]<=26'd11160234; ROM3[7746]<=26'd9771670; ROM4[7746]<=26'd23496175;
ROM1[7747]<=26'd2058151; ROM2[7747]<=26'd11162613; ROM3[7747]<=26'd9768741; ROM4[7747]<=26'd23497218;
ROM1[7748]<=26'd2072997; ROM2[7748]<=26'd11167149; ROM3[7748]<=26'd9768033; ROM4[7748]<=26'd23498614;
ROM1[7749]<=26'd2071748; ROM2[7749]<=26'd11167488; ROM3[7749]<=26'd9766543; ROM4[7749]<=26'd23497301;
ROM1[7750]<=26'd2059399; ROM2[7750]<=26'd11162226; ROM3[7750]<=26'd9762523; ROM4[7750]<=26'd23492247;
ROM1[7751]<=26'd2053036; ROM2[7751]<=26'd11163683; ROM3[7751]<=26'd9766275; ROM4[7751]<=26'd23492514;
ROM1[7752]<=26'd2049199; ROM2[7752]<=26'd11163695; ROM3[7752]<=26'd9770120; ROM4[7752]<=26'd23495114;
ROM1[7753]<=26'd2043434; ROM2[7753]<=26'd11160894; ROM3[7753]<=26'd9773073; ROM4[7753]<=26'd23495933;
ROM1[7754]<=26'd2042069; ROM2[7754]<=26'd11162839; ROM3[7754]<=26'd9775887; ROM4[7754]<=26'd23497938;
ROM1[7755]<=26'd2047650; ROM2[7755]<=26'd11164514; ROM3[7755]<=26'd9774501; ROM4[7755]<=26'd23497283;
ROM1[7756]<=26'd2059631; ROM2[7756]<=26'd11164652; ROM3[7756]<=26'd9768582; ROM4[7756]<=26'd23497256;
ROM1[7757]<=26'd2070802; ROM2[7757]<=26'd11170990; ROM3[7757]<=26'd9770593; ROM4[7757]<=26'd23503086;
ROM1[7758]<=26'd2069306; ROM2[7758]<=26'd11174356; ROM3[7758]<=26'd9776769; ROM4[7758]<=26'd23505637;
ROM1[7759]<=26'd2051154; ROM2[7759]<=26'd11162086; ROM3[7759]<=26'd9769272; ROM4[7759]<=26'd23496494;
ROM1[7760]<=26'd2033166; ROM2[7760]<=26'd11151591; ROM3[7760]<=26'd9761962; ROM4[7760]<=26'd23487122;
ROM1[7761]<=26'd2021434; ROM2[7761]<=26'd11145585; ROM3[7761]<=26'd9759262; ROM4[7761]<=26'd23480365;
ROM1[7762]<=26'd2018142; ROM2[7762]<=26'd11143537; ROM3[7762]<=26'd9757637; ROM4[7762]<=26'd23478440;
ROM1[7763]<=26'd2026145; ROM2[7763]<=26'd11148066; ROM3[7763]<=26'd9757816; ROM4[7763]<=26'd23481621;
ROM1[7764]<=26'd2037872; ROM2[7764]<=26'd11150633; ROM3[7764]<=26'd9753782; ROM4[7764]<=26'd23480355;
ROM1[7765]<=26'd2045210; ROM2[7765]<=26'd11151652; ROM3[7765]<=26'd9748348; ROM4[7765]<=26'd23479254;
ROM1[7766]<=26'd2040747; ROM2[7766]<=26'd11151326; ROM3[7766]<=26'd9747274; ROM4[7766]<=26'd23478579;
ROM1[7767]<=26'd2032920; ROM2[7767]<=26'd11152829; ROM3[7767]<=26'd9751203; ROM4[7767]<=26'd23479400;
ROM1[7768]<=26'd2024820; ROM2[7768]<=26'd11150841; ROM3[7768]<=26'd9751880; ROM4[7768]<=26'd23477187;
ROM1[7769]<=26'd2018882; ROM2[7769]<=26'd11148906; ROM3[7769]<=26'd9752274; ROM4[7769]<=26'd23475568;
ROM1[7770]<=26'd2012366; ROM2[7770]<=26'd11146843; ROM3[7770]<=26'd9753455; ROM4[7770]<=26'd23474645;
ROM1[7771]<=26'd2009225; ROM2[7771]<=26'd11142301; ROM3[7771]<=26'd9749973; ROM4[7771]<=26'd23470621;
ROM1[7772]<=26'd2021706; ROM2[7772]<=26'd11146398; ROM3[7772]<=26'd9748856; ROM4[7772]<=26'd23471705;
ROM1[7773]<=26'd2038632; ROM2[7773]<=26'd11151969; ROM3[7773]<=26'd9747483; ROM4[7773]<=26'd23476472;
ROM1[7774]<=26'd2033012; ROM2[7774]<=26'd11145895; ROM3[7774]<=26'd9740812; ROM4[7774]<=26'd23471002;
ROM1[7775]<=26'd2020179; ROM2[7775]<=26'd11139050; ROM3[7775]<=26'd9737391; ROM4[7775]<=26'd23463408;
ROM1[7776]<=26'd2014079; ROM2[7776]<=26'd11138429; ROM3[7776]<=26'd9742477; ROM4[7776]<=26'd23465365;
ROM1[7777]<=26'd2010046; ROM2[7777]<=26'd11140832; ROM3[7777]<=26'd9746393; ROM4[7777]<=26'd23467819;
ROM1[7778]<=26'd2005746; ROM2[7778]<=26'd11142258; ROM3[7778]<=26'd9748560; ROM4[7778]<=26'd23468610;
ROM1[7779]<=26'd2006628; ROM2[7779]<=26'd11142637; ROM3[7779]<=26'd9749465; ROM4[7779]<=26'd23469581;
ROM1[7780]<=26'd2015672; ROM2[7780]<=26'd11147043; ROM3[7780]<=26'd9749745; ROM4[7780]<=26'd23473612;
ROM1[7781]<=26'd2027372; ROM2[7781]<=26'd11148848; ROM3[7781]<=26'd9746705; ROM4[7781]<=26'd23474165;
ROM1[7782]<=26'd2039328; ROM2[7782]<=26'd11155589; ROM3[7782]<=26'd9751052; ROM4[7782]<=26'd23480342;
ROM1[7783]<=26'd2041858; ROM2[7783]<=26'd11163482; ROM3[7783]<=26'd9758867; ROM4[7783]<=26'd23489165;
ROM1[7784]<=26'd2024844; ROM2[7784]<=26'd11151941; ROM3[7784]<=26'd9750198; ROM4[7784]<=26'd23478872;
ROM1[7785]<=26'd2009666; ROM2[7785]<=26'd11141212; ROM3[7785]<=26'd9743676; ROM4[7785]<=26'd23468752;
ROM1[7786]<=26'd2001287; ROM2[7786]<=26'd11138246; ROM3[7786]<=26'd9743734; ROM4[7786]<=26'd23465485;
ROM1[7787]<=26'd1995752; ROM2[7787]<=26'd11135119; ROM3[7787]<=26'd9742609; ROM4[7787]<=26'd23462029;
ROM1[7788]<=26'd2000688; ROM2[7788]<=26'd11137822; ROM3[7788]<=26'd9743326; ROM4[7788]<=26'd23464000;
ROM1[7789]<=26'd2017073; ROM2[7789]<=26'd11143177; ROM3[7789]<=26'd9743659; ROM4[7789]<=26'd23468379;
ROM1[7790]<=26'd2030903; ROM2[7790]<=26'd11145140; ROM3[7790]<=26'd9742545; ROM4[7790]<=26'd23471136;
ROM1[7791]<=26'd2025885; ROM2[7791]<=26'd11143062; ROM3[7791]<=26'd9745334; ROM4[7791]<=26'd23470459;
ROM1[7792]<=26'd2015432; ROM2[7792]<=26'd11141129; ROM3[7792]<=26'd9749613; ROM4[7792]<=26'd23469752;
ROM1[7793]<=26'd2007012; ROM2[7793]<=26'd11138491; ROM3[7793]<=26'd9752644; ROM4[7793]<=26'd23469049;
ROM1[7794]<=26'd2004223; ROM2[7794]<=26'd11140972; ROM3[7794]<=26'd9759054; ROM4[7794]<=26'd23472907;
ROM1[7795]<=26'd2005113; ROM2[7795]<=26'd11144355; ROM3[7795]<=26'd9765456; ROM4[7795]<=26'd23478021;
ROM1[7796]<=26'd2008739; ROM2[7796]<=26'd11145680; ROM3[7796]<=26'd9767367; ROM4[7796]<=26'd23480073;
ROM1[7797]<=26'd2016409; ROM2[7797]<=26'd11146345; ROM3[7797]<=26'd9762589; ROM4[7797]<=26'd23479840;
ROM1[7798]<=26'd2026603; ROM2[7798]<=26'd11144926; ROM3[7798]<=26'd9756560; ROM4[7798]<=26'd23479494;
ROM1[7799]<=26'd2026433; ROM2[7799]<=26'd11143870; ROM3[7799]<=26'd9753422; ROM4[7799]<=26'd23478560;
ROM1[7800]<=26'd2024590; ROM2[7800]<=26'd11148759; ROM3[7800]<=26'd9758432; ROM4[7800]<=26'd23482117;
ROM1[7801]<=26'd2022418; ROM2[7801]<=26'd11152473; ROM3[7801]<=26'd9766352; ROM4[7801]<=26'd23486979;
ROM1[7802]<=26'd2021541; ROM2[7802]<=26'd11157006; ROM3[7802]<=26'd9773135; ROM4[7802]<=26'd23492148;
ROM1[7803]<=26'd2009752; ROM2[7803]<=26'd11149191; ROM3[7803]<=26'd9768500; ROM4[7803]<=26'd23485477;
ROM1[7804]<=26'd2004185; ROM2[7804]<=26'd11142064; ROM3[7804]<=26'd9764535; ROM4[7804]<=26'd23478950;
ROM1[7805]<=26'd2018360; ROM2[7805]<=26'd11150350; ROM3[7805]<=26'd9769080; ROM4[7805]<=26'd23485365;
ROM1[7806]<=26'd2023573; ROM2[7806]<=26'd11144795; ROM3[7806]<=26'd9755581; ROM4[7806]<=26'd23477817;
ROM1[7807]<=26'd2027028; ROM2[7807]<=26'd11143108; ROM3[7807]<=26'd9750653; ROM4[7807]<=26'd23475728;
ROM1[7808]<=26'd2024649; ROM2[7808]<=26'd11147185; ROM3[7808]<=26'd9756724; ROM4[7808]<=26'd23480013;
ROM1[7809]<=26'd2014385; ROM2[7809]<=26'd11143383; ROM3[7809]<=26'd9758216; ROM4[7809]<=26'd23478089;
ROM1[7810]<=26'd2003492; ROM2[7810]<=26'd11137321; ROM3[7810]<=26'd9755142; ROM4[7810]<=26'd23471809;
ROM1[7811]<=26'd1996076; ROM2[7811]<=26'd11135266; ROM3[7811]<=26'd9753392; ROM4[7811]<=26'd23470254;
ROM1[7812]<=26'd1994753; ROM2[7812]<=26'd11133043; ROM3[7812]<=26'd9752868; ROM4[7812]<=26'd23469751;
ROM1[7813]<=26'd1994688; ROM2[7813]<=26'd11130392; ROM3[7813]<=26'd9745074; ROM4[7813]<=26'd23463155;
ROM1[7814]<=26'd2008065; ROM2[7814]<=26'd11135730; ROM3[7814]<=26'd9742440; ROM4[7814]<=26'd23465904;
ROM1[7815]<=26'd2022333; ROM2[7815]<=26'd11141071; ROM3[7815]<=26'd9743056; ROM4[7815]<=26'd23470411;
ROM1[7816]<=26'd2015061; ROM2[7816]<=26'd11137899; ROM3[7816]<=26'd9738064; ROM4[7816]<=26'd23466340;
ROM1[7817]<=26'd2005146; ROM2[7817]<=26'd11135593; ROM3[7817]<=26'd9737749; ROM4[7817]<=26'd23462701;
ROM1[7818]<=26'd2005766; ROM2[7818]<=26'd11141823; ROM3[7818]<=26'd9750028; ROM4[7818]<=26'd23470270;
ROM1[7819]<=26'd2001665; ROM2[7819]<=26'd11145902; ROM3[7819]<=26'd9757373; ROM4[7819]<=26'd23475741;
ROM1[7820]<=26'd1992804; ROM2[7820]<=26'd11140947; ROM3[7820]<=26'd9752030; ROM4[7820]<=26'd23470459;
ROM1[7821]<=26'd1990106; ROM2[7821]<=26'd11134906; ROM3[7821]<=26'd9748036; ROM4[7821]<=26'd23466177;
ROM1[7822]<=26'd1997436; ROM2[7822]<=26'd11132318; ROM3[7822]<=26'd9744005; ROM4[7822]<=26'd23463506;
ROM1[7823]<=26'd2013257; ROM2[7823]<=26'd11135753; ROM3[7823]<=26'd9739511; ROM4[7823]<=26'd23464569;
ROM1[7824]<=26'd2021017; ROM2[7824]<=26'd11143797; ROM3[7824]<=26'd9746263; ROM4[7824]<=26'd23472026;
ROM1[7825]<=26'd2016374; ROM2[7825]<=26'd11145622; ROM3[7825]<=26'd9751035; ROM4[7825]<=26'd23476341;
ROM1[7826]<=26'd2008411; ROM2[7826]<=26'd11141880; ROM3[7826]<=26'd9750645; ROM4[7826]<=26'd23473399;
ROM1[7827]<=26'd2001227; ROM2[7827]<=26'd11140355; ROM3[7827]<=26'd9750015; ROM4[7827]<=26'd23469896;
ROM1[7828]<=26'd2001994; ROM2[7828]<=26'd11148878; ROM3[7828]<=26'd9759729; ROM4[7828]<=26'd23478886;
ROM1[7829]<=26'd2010350; ROM2[7829]<=26'd11156142; ROM3[7829]<=26'd9768672; ROM4[7829]<=26'd23487803;
ROM1[7830]<=26'd2002062; ROM2[7830]<=26'd11142917; ROM3[7830]<=26'd9751902; ROM4[7830]<=26'd23473204;
ROM1[7831]<=26'd2002634; ROM2[7831]<=26'd11134218; ROM3[7831]<=26'd9737458; ROM4[7831]<=26'd23463535;
ROM1[7832]<=26'd2005468; ROM2[7832]<=26'd11131477; ROM3[7832]<=26'd9733300; ROM4[7832]<=26'd23461643;
ROM1[7833]<=26'd1997108; ROM2[7833]<=26'd11128829; ROM3[7833]<=26'd9730372; ROM4[7833]<=26'd23457085;
ROM1[7834]<=26'd1995473; ROM2[7834]<=26'd11136875; ROM3[7834]<=26'd9739777; ROM4[7834]<=26'd23464320;
ROM1[7835]<=26'd1995360; ROM2[7835]<=26'd11140365; ROM3[7835]<=26'd9747227; ROM4[7835]<=26'd23468834;
ROM1[7836]<=26'd1983704; ROM2[7836]<=26'd11131980; ROM3[7836]<=26'd9741830; ROM4[7836]<=26'd23461205;
ROM1[7837]<=26'd1975969; ROM2[7837]<=26'd11126319; ROM3[7837]<=26'd9736788; ROM4[7837]<=26'd23455600;
ROM1[7838]<=26'd1986160; ROM2[7838]<=26'd11131906; ROM3[7838]<=26'd9740905; ROM4[7838]<=26'd23461080;
ROM1[7839]<=26'd2002309; ROM2[7839]<=26'd11138694; ROM3[7839]<=26'd9742460; ROM4[7839]<=26'd23467133;
ROM1[7840]<=26'd2011312; ROM2[7840]<=26'd11141057; ROM3[7840]<=26'd9738991; ROM4[7840]<=26'd23468218;
ROM1[7841]<=26'd2007149; ROM2[7841]<=26'd11140510; ROM3[7841]<=26'd9740027; ROM4[7841]<=26'd23470325;
ROM1[7842]<=26'd2003645; ROM2[7842]<=26'd11143417; ROM3[7842]<=26'd9746935; ROM4[7842]<=26'd23475054;
ROM1[7843]<=26'd1998683; ROM2[7843]<=26'd11142834; ROM3[7843]<=26'd9749720; ROM4[7843]<=26'd23473829;
ROM1[7844]<=26'd1985939; ROM2[7844]<=26'd11134295; ROM3[7844]<=26'd9744549; ROM4[7844]<=26'd23465941;
ROM1[7845]<=26'd1973739; ROM2[7845]<=26'd11127538; ROM3[7845]<=26'd9740587; ROM4[7845]<=26'd23458478;
ROM1[7846]<=26'd1975241; ROM2[7846]<=26'd11128074; ROM3[7846]<=26'd9739659; ROM4[7846]<=26'd23459253;
ROM1[7847]<=26'd1985133; ROM2[7847]<=26'd11128543; ROM3[7847]<=26'd9736751; ROM4[7847]<=26'd23460685;
ROM1[7848]<=26'd1999651; ROM2[7848]<=26'd11131610; ROM3[7848]<=26'd9735496; ROM4[7848]<=26'd23462861;
ROM1[7849]<=26'd2007734; ROM2[7849]<=26'd11137627; ROM3[7849]<=26'd9740002; ROM4[7849]<=26'd23467309;
ROM1[7850]<=26'd2004504; ROM2[7850]<=26'd11140969; ROM3[7850]<=26'd9744710; ROM4[7850]<=26'd23469155;
ROM1[7851]<=26'd1996457; ROM2[7851]<=26'd11140105; ROM3[7851]<=26'd9747670; ROM4[7851]<=26'd23468003;
ROM1[7852]<=26'd1988198; ROM2[7852]<=26'd11136199; ROM3[7852]<=26'd9747789; ROM4[7852]<=26'd23465976;
ROM1[7853]<=26'd1983763; ROM2[7853]<=26'd11134646; ROM3[7853]<=26'd9750309; ROM4[7853]<=26'd23467224;
ROM1[7854]<=26'd1984075; ROM2[7854]<=26'd11133805; ROM3[7854]<=26'd9751013; ROM4[7854]<=26'd23466608;
ROM1[7855]<=26'd1991789; ROM2[7855]<=26'd11135710; ROM3[7855]<=26'd9750989; ROM4[7855]<=26'd23467399;
ROM1[7856]<=26'd2006513; ROM2[7856]<=26'd11138463; ROM3[7856]<=26'd9748124; ROM4[7856]<=26'd23468601;
ROM1[7857]<=26'd2008528; ROM2[7857]<=26'd11138045; ROM3[7857]<=26'd9741595; ROM4[7857]<=26'd23466701;
ROM1[7858]<=26'd1999970; ROM2[7858]<=26'd11134684; ROM3[7858]<=26'd9740002; ROM4[7858]<=26'd23463568;
ROM1[7859]<=26'd1990870; ROM2[7859]<=26'd11131409; ROM3[7859]<=26'd9740535; ROM4[7859]<=26'd23462289;
ROM1[7860]<=26'd1987308; ROM2[7860]<=26'd11133689; ROM3[7860]<=26'd9744957; ROM4[7860]<=26'd23465163;
ROM1[7861]<=26'd1983029; ROM2[7861]<=26'd11136025; ROM3[7861]<=26'd9751898; ROM4[7861]<=26'd23467862;
ROM1[7862]<=26'd1976860; ROM2[7862]<=26'd11133517; ROM3[7862]<=26'd9750612; ROM4[7862]<=26'd23466096;
ROM1[7863]<=26'd1975313; ROM2[7863]<=26'd11129772; ROM3[7863]<=26'd9744225; ROM4[7863]<=26'd23460960;
ROM1[7864]<=26'd1988112; ROM2[7864]<=26'd11132794; ROM3[7864]<=26'd9742057; ROM4[7864]<=26'd23460602;
ROM1[7865]<=26'd1996060; ROM2[7865]<=26'd11131999; ROM3[7865]<=26'd9735530; ROM4[7865]<=26'd23458514;
ROM1[7866]<=26'd1987851; ROM2[7866]<=26'd11126622; ROM3[7866]<=26'd9730365; ROM4[7866]<=26'd23453320;
ROM1[7867]<=26'd1982723; ROM2[7867]<=26'd11127365; ROM3[7867]<=26'd9734074; ROM4[7867]<=26'd23454065;
ROM1[7868]<=26'd1983781; ROM2[7868]<=26'd11134116; ROM3[7868]<=26'd9742633; ROM4[7868]<=26'd23460344;
ROM1[7869]<=26'd1981329; ROM2[7869]<=26'd11135345; ROM3[7869]<=26'd9745039; ROM4[7869]<=26'd23461777;
ROM1[7870]<=26'd1974474; ROM2[7870]<=26'd11130897; ROM3[7870]<=26'd9742244; ROM4[7870]<=26'd23458423;
ROM1[7871]<=26'd1976317; ROM2[7871]<=26'd11131199; ROM3[7871]<=26'd9743069; ROM4[7871]<=26'd23459008;
ROM1[7872]<=26'd1981925; ROM2[7872]<=26'd11126974; ROM3[7872]<=26'd9733781; ROM4[7872]<=26'd23453320;
ROM1[7873]<=26'd1992102; ROM2[7873]<=26'd11126296; ROM3[7873]<=26'd9725341; ROM4[7873]<=26'd23450648;
ROM1[7874]<=26'd1994135; ROM2[7874]<=26'd11129091; ROM3[7874]<=26'd9725935; ROM4[7874]<=26'd23452447;
ROM1[7875]<=26'd1986535; ROM2[7875]<=26'd11129663; ROM3[7875]<=26'd9726976; ROM4[7875]<=26'd23451641;
ROM1[7876]<=26'd1975658; ROM2[7876]<=26'd11125878; ROM3[7876]<=26'd9728152; ROM4[7876]<=26'd23450661;
ROM1[7877]<=26'd1971156; ROM2[7877]<=26'd11125246; ROM3[7877]<=26'd9731337; ROM4[7877]<=26'd23451057;
ROM1[7878]<=26'd1969168; ROM2[7878]<=26'd11129362; ROM3[7878]<=26'd9735692; ROM4[7878]<=26'd23453614;
ROM1[7879]<=26'd1970555; ROM2[7879]<=26'd11132467; ROM3[7879]<=26'd9736996; ROM4[7879]<=26'd23455757;
ROM1[7880]<=26'd1978760; ROM2[7880]<=26'd11136841; ROM3[7880]<=26'd9736255; ROM4[7880]<=26'd23457826;
ROM1[7881]<=26'd1989196; ROM2[7881]<=26'd11137398; ROM3[7881]<=26'd9732630; ROM4[7881]<=26'd23457554;
ROM1[7882]<=26'd1992103; ROM2[7882]<=26'd11133584; ROM3[7882]<=26'd9729464; ROM4[7882]<=26'd23456254;
ROM1[7883]<=26'd1989347; ROM2[7883]<=26'd11132760; ROM3[7883]<=26'd9731999; ROM4[7883]<=26'd23457685;
ROM1[7884]<=26'd1985025; ROM2[7884]<=26'd11135248; ROM3[7884]<=26'd9737757; ROM4[7884]<=26'd23460507;
ROM1[7885]<=26'd1989212; ROM2[7885]<=26'd11142132; ROM3[7885]<=26'd9751124; ROM4[7885]<=26'd23468098;
ROM1[7886]<=26'd1983799; ROM2[7886]<=26'd11140590; ROM3[7886]<=26'd9753945; ROM4[7886]<=26'd23467164;
ROM1[7887]<=26'd1963796; ROM2[7887]<=26'd11123698; ROM3[7887]<=26'd9737821; ROM4[7887]<=26'd23451042;
ROM1[7888]<=26'd1967646; ROM2[7888]<=26'd11121839; ROM3[7888]<=26'd9733267; ROM4[7888]<=26'd23447998;
ROM1[7889]<=26'd1979841; ROM2[7889]<=26'd11123916; ROM3[7889]<=26'd9727507; ROM4[7889]<=26'd23448664;
ROM1[7890]<=26'd1984428; ROM2[7890]<=26'd11121326; ROM3[7890]<=26'd9719230; ROM4[7890]<=26'd23445213;
ROM1[7891]<=26'd1986574; ROM2[7891]<=26'd11124863; ROM3[7891]<=26'd9721730; ROM4[7891]<=26'd23448982;
ROM1[7892]<=26'd1979167; ROM2[7892]<=26'd11123682; ROM3[7892]<=26'd9723573; ROM4[7892]<=26'd23449743;
ROM1[7893]<=26'd1967787; ROM2[7893]<=26'd11118575; ROM3[7893]<=26'd9723751; ROM4[7893]<=26'd23445883;
ROM1[7894]<=26'd1966503; ROM2[7894]<=26'd11121866; ROM3[7894]<=26'd9731044; ROM4[7894]<=26'd23450069;
ROM1[7895]<=26'd1971710; ROM2[7895]<=26'd11130161; ROM3[7895]<=26'd9741707; ROM4[7895]<=26'd23457464;
ROM1[7896]<=26'd1974707; ROM2[7896]<=26'd11133437; ROM3[7896]<=26'd9743853; ROM4[7896]<=26'd23460128;
ROM1[7897]<=26'd1977772; ROM2[7897]<=26'd11127825; ROM3[7897]<=26'd9731153; ROM4[7897]<=26'd23453808;
ROM1[7898]<=26'd1983158; ROM2[7898]<=26'd11121431; ROM3[7898]<=26'd9716412; ROM4[7898]<=26'd23445104;
ROM1[7899]<=26'd1984934; ROM2[7899]<=26'd11123835; ROM3[7899]<=26'd9718635; ROM4[7899]<=26'd23448320;
ROM1[7900]<=26'd1976154; ROM2[7900]<=26'd11120814; ROM3[7900]<=26'd9720116; ROM4[7900]<=26'd23447611;
ROM1[7901]<=26'd1966849; ROM2[7901]<=26'd11117431; ROM3[7901]<=26'd9722534; ROM4[7901]<=26'd23446342;
ROM1[7902]<=26'd1966764; ROM2[7902]<=26'd11123664; ROM3[7902]<=26'd9731952; ROM4[7902]<=26'd23452890;
ROM1[7903]<=26'd1962407; ROM2[7903]<=26'd11122676; ROM3[7903]<=26'd9735940; ROM4[7903]<=26'd23454133;
ROM1[7904]<=26'd1960135; ROM2[7904]<=26'd11118998; ROM3[7904]<=26'd9732580; ROM4[7904]<=26'd23451107;
ROM1[7905]<=26'd1971225; ROM2[7905]<=26'd11124591; ROM3[7905]<=26'd9733604; ROM4[7905]<=26'd23455058;
ROM1[7906]<=26'd1986142; ROM2[7906]<=26'd11128209; ROM3[7906]<=26'd9732782; ROM4[7906]<=26'd23457382;
ROM1[7907]<=26'd1988534; ROM2[7907]<=26'd11126767; ROM3[7907]<=26'd9728214; ROM4[7907]<=26'd23455378;
ROM1[7908]<=26'd1987051; ROM2[7908]<=26'd11129392; ROM3[7908]<=26'd9733313; ROM4[7908]<=26'd23459493;
ROM1[7909]<=26'd1984428; ROM2[7909]<=26'd11133062; ROM3[7909]<=26'd9741323; ROM4[7909]<=26'd23463204;
ROM1[7910]<=26'd1981166; ROM2[7910]<=26'd11134055; ROM3[7910]<=26'd9744606; ROM4[7910]<=26'd23465136;
ROM1[7911]<=26'd1977613; ROM2[7911]<=26'd11134657; ROM3[7911]<=26'd9747283; ROM4[7911]<=26'd23466734;
ROM1[7912]<=26'd1973833; ROM2[7912]<=26'd11133388; ROM3[7912]<=26'd9746212; ROM4[7912]<=26'd23464636;
ROM1[7913]<=26'd1975089; ROM2[7913]<=26'd11131098; ROM3[7913]<=26'd9741388; ROM4[7913]<=26'd23461752;
ROM1[7914]<=26'd1989541; ROM2[7914]<=26'd11134879; ROM3[7914]<=26'd9740366; ROM4[7914]<=26'd23463839;
ROM1[7915]<=26'd2007698; ROM2[7915]<=26'd11143601; ROM3[7915]<=26'd9745249; ROM4[7915]<=26'd23471685;
ROM1[7916]<=26'd2005639; ROM2[7916]<=26'd11141994; ROM3[7916]<=26'd9744618; ROM4[7916]<=26'd23471156;
ROM1[7917]<=26'd1993850; ROM2[7917]<=26'd11135708; ROM3[7917]<=26'd9740680; ROM4[7917]<=26'd23467317;
ROM1[7918]<=26'd1983228; ROM2[7918]<=26'd11131185; ROM3[7918]<=26'd9739220; ROM4[7918]<=26'd23464923;
ROM1[7919]<=26'd1972599; ROM2[7919]<=26'd11123922; ROM3[7919]<=26'd9737362; ROM4[7919]<=26'd23459971;
ROM1[7920]<=26'd1971884; ROM2[7920]<=26'd11126560; ROM3[7920]<=26'd9744252; ROM4[7920]<=26'd23462688;
ROM1[7921]<=26'd1973147; ROM2[7921]<=26'd11126206; ROM3[7921]<=26'd9742474; ROM4[7921]<=26'd23460659;
ROM1[7922]<=26'd1981338; ROM2[7922]<=26'd11124965; ROM3[7922]<=26'd9735515; ROM4[7922]<=26'd23457627;
ROM1[7923]<=26'd1993548; ROM2[7923]<=26'd11128391; ROM3[7923]<=26'd9730072; ROM4[7923]<=26'd23457512;
ROM1[7924]<=26'd1991911; ROM2[7924]<=26'd11128237; ROM3[7924]<=26'd9728773; ROM4[7924]<=26'd23457015;
ROM1[7925]<=26'd1990203; ROM2[7925]<=26'd11132208; ROM3[7925]<=26'd9736285; ROM4[7925]<=26'd23461324;
ROM1[7926]<=26'd1987688; ROM2[7926]<=26'd11135135; ROM3[7926]<=26'd9745155; ROM4[7926]<=26'd23466661;
ROM1[7927]<=26'd1983554; ROM2[7927]<=26'd11134206; ROM3[7927]<=26'd9747959; ROM4[7927]<=26'd23466407;
ROM1[7928]<=26'd1975673; ROM2[7928]<=26'd11131933; ROM3[7928]<=26'd9746652; ROM4[7928]<=26'd23461899;
ROM1[7929]<=26'd1973284; ROM2[7929]<=26'd11130504; ROM3[7929]<=26'd9745289; ROM4[7929]<=26'd23460327;
ROM1[7930]<=26'd1984627; ROM2[7930]<=26'd11134229; ROM3[7930]<=26'd9744074; ROM4[7930]<=26'd23462318;
ROM1[7931]<=26'd1996970; ROM2[7931]<=26'd11135719; ROM3[7931]<=26'd9737894; ROM4[7931]<=26'd23460576;
ROM1[7932]<=26'd1998123; ROM2[7932]<=26'd11131932; ROM3[7932]<=26'd9730187; ROM4[7932]<=26'd23456902;
ROM1[7933]<=26'd1996865; ROM2[7933]<=26'd11135581; ROM3[7933]<=26'd9733449; ROM4[7933]<=26'd23459931;
ROM1[7934]<=26'd1993400; ROM2[7934]<=26'd11140286; ROM3[7934]<=26'd9739040; ROM4[7934]<=26'd23462746;
ROM1[7935]<=26'd1982151; ROM2[7935]<=26'd11136500; ROM3[7935]<=26'd9737525; ROM4[7935]<=26'd23458709;
ROM1[7936]<=26'd1969719; ROM2[7936]<=26'd11129962; ROM3[7936]<=26'd9734035; ROM4[7936]<=26'd23453463;
ROM1[7937]<=26'd1971898; ROM2[7937]<=26'd11134116; ROM3[7937]<=26'd9738383; ROM4[7937]<=26'd23456926;
ROM1[7938]<=26'd1974278; ROM2[7938]<=26'd11133363; ROM3[7938]<=26'd9736640; ROM4[7938]<=26'd23455789;
ROM1[7939]<=26'd1978760; ROM2[7939]<=26'd11127897; ROM3[7939]<=26'd9725926; ROM4[7939]<=26'd23449610;
ROM1[7940]<=26'd1992083; ROM2[7940]<=26'd11132172; ROM3[7940]<=26'd9725108; ROM4[7940]<=26'd23451331;
ROM1[7941]<=26'd1988807; ROM2[7941]<=26'd11130651; ROM3[7941]<=26'd9727191; ROM4[7941]<=26'd23452002;
ROM1[7942]<=26'd1981777; ROM2[7942]<=26'd11129981; ROM3[7942]<=26'd9728357; ROM4[7942]<=26'd23450776;
ROM1[7943]<=26'd1979151; ROM2[7943]<=26'd11132751; ROM3[7943]<=26'd9734954; ROM4[7943]<=26'd23453417;
ROM1[7944]<=26'd1974185; ROM2[7944]<=26'd11133525; ROM3[7944]<=26'd9738601; ROM4[7944]<=26'd23455950;
ROM1[7945]<=26'd1967789; ROM2[7945]<=26'd11129632; ROM3[7945]<=26'd9737504; ROM4[7945]<=26'd23451326;
ROM1[7946]<=26'd1966909; ROM2[7946]<=26'd11123623; ROM3[7946]<=26'd9734609; ROM4[7946]<=26'd23447233;
ROM1[7947]<=26'd1978870; ROM2[7947]<=26'd11127858; ROM3[7947]<=26'd9732484; ROM4[7947]<=26'd23449207;
ROM1[7948]<=26'd1994032; ROM2[7948]<=26'd11132930; ROM3[7948]<=26'd9730491; ROM4[7948]<=26'd23451059;
ROM1[7949]<=26'd1995525; ROM2[7949]<=26'd11132102; ROM3[7949]<=26'd9727749; ROM4[7949]<=26'd23451613;
ROM1[7950]<=26'd1987846; ROM2[7950]<=26'd11131254; ROM3[7950]<=26'd9728582; ROM4[7950]<=26'd23452254;
ROM1[7951]<=26'd1987696; ROM2[7951]<=26'd11137738; ROM3[7951]<=26'd9737921; ROM4[7951]<=26'd23459558;
ROM1[7952]<=26'd1986779; ROM2[7952]<=26'd11141872; ROM3[7952]<=26'd9744397; ROM4[7952]<=26'd23464675;
ROM1[7953]<=26'd1969852; ROM2[7953]<=26'd11131225; ROM3[7953]<=26'd9736723; ROM4[7953]<=26'd23455781;
ROM1[7954]<=26'd1965219; ROM2[7954]<=26'd11127126; ROM3[7954]<=26'd9733315; ROM4[7954]<=26'd23452254;
ROM1[7955]<=26'd1974035; ROM2[7955]<=26'd11127333; ROM3[7955]<=26'd9731813; ROM4[7955]<=26'd23452249;
ROM1[7956]<=26'd1988395; ROM2[7956]<=26'd11128351; ROM3[7956]<=26'd9725485; ROM4[7956]<=26'd23451816;
ROM1[7957]<=26'd1999903; ROM2[7957]<=26'd11135515; ROM3[7957]<=26'd9728666; ROM4[7957]<=26'd23457987;
ROM1[7958]<=26'd1997394; ROM2[7958]<=26'd11139270; ROM3[7958]<=26'd9733589; ROM4[7958]<=26'd23462560;
ROM1[7959]<=26'd1987912; ROM2[7959]<=26'd11136445; ROM3[7959]<=26'd9734165; ROM4[7959]<=26'd23461433;
ROM1[7960]<=26'd1979014; ROM2[7960]<=26'd11131617; ROM3[7960]<=26'd9734792; ROM4[7960]<=26'd23458974;
ROM1[7961]<=26'd1974778; ROM2[7961]<=26'd11131816; ROM3[7961]<=26'd9740357; ROM4[7961]<=26'd23460646;
ROM1[7962]<=26'd1976463; ROM2[7962]<=26'd11133164; ROM3[7962]<=26'd9742977; ROM4[7962]<=26'd23463165;
ROM1[7963]<=26'd1983925; ROM2[7963]<=26'd11136458; ROM3[7963]<=26'd9741674; ROM4[7963]<=26'd23465942;
ROM1[7964]<=26'd1997313; ROM2[7964]<=26'd11139210; ROM3[7964]<=26'd9738727; ROM4[7964]<=26'd23467122;
ROM1[7965]<=26'd2002386; ROM2[7965]<=26'd11136900; ROM3[7965]<=26'd9730125; ROM4[7965]<=26'd23462526;
ROM1[7966]<=26'd1995691; ROM2[7966]<=26'd11133648; ROM3[7966]<=26'd9727714; ROM4[7966]<=26'd23458421;
ROM1[7967]<=26'd1987435; ROM2[7967]<=26'd11132518; ROM3[7967]<=26'd9732878; ROM4[7967]<=26'd23459179;
ROM1[7968]<=26'd1975908; ROM2[7968]<=26'd11128474; ROM3[7968]<=26'd9732866; ROM4[7968]<=26'd23456888;
ROM1[7969]<=26'd1973264; ROM2[7969]<=26'd11131286; ROM3[7969]<=26'd9738240; ROM4[7969]<=26'd23460342;
ROM1[7970]<=26'd1970892; ROM2[7970]<=26'd11132462; ROM3[7970]<=26'd9741708; ROM4[7970]<=26'd23460884;
ROM1[7971]<=26'd1970153; ROM2[7971]<=26'd11129716; ROM3[7971]<=26'd9737199; ROM4[7971]<=26'd23457775;
ROM1[7972]<=26'd1981779; ROM2[7972]<=26'd11130688; ROM3[7972]<=26'd9734776; ROM4[7972]<=26'd23458253;
ROM1[7973]<=26'd1992254; ROM2[7973]<=26'd11131533; ROM3[7973]<=26'd9729519; ROM4[7973]<=26'd23459472;
ROM1[7974]<=26'd1989209; ROM2[7974]<=26'd11128400; ROM3[7974]<=26'd9724753; ROM4[7974]<=26'd23457056;
ROM1[7975]<=26'd1983248; ROM2[7975]<=26'd11128395; ROM3[7975]<=26'd9727440; ROM4[7975]<=26'd23457451;
ROM1[7976]<=26'd1978358; ROM2[7976]<=26'd11129351; ROM3[7976]<=26'd9733144; ROM4[7976]<=26'd23460164;
ROM1[7977]<=26'd1973463; ROM2[7977]<=26'd11127440; ROM3[7977]<=26'd9733826; ROM4[7977]<=26'd23458389;
ROM1[7978]<=26'd1970816; ROM2[7978]<=26'd11130133; ROM3[7978]<=26'd9739364; ROM4[7978]<=26'd23461816;
ROM1[7979]<=26'd1974343; ROM2[7979]<=26'd11133880; ROM3[7979]<=26'd9743793; ROM4[7979]<=26'd23465619;
ROM1[7980]<=26'd1993401; ROM2[7980]<=26'd11146929; ROM3[7980]<=26'd9751139; ROM4[7980]<=26'd23475408;
ROM1[7981]<=26'd2001416; ROM2[7981]<=26'd11144643; ROM3[7981]<=26'd9743076; ROM4[7981]<=26'd23469859;
ROM1[7982]<=26'd1990196; ROM2[7982]<=26'd11129109; ROM3[7982]<=26'd9724088; ROM4[7982]<=26'd23453229;
ROM1[7983]<=26'd1982428; ROM2[7983]<=26'd11127466; ROM3[7983]<=26'd9722545; ROM4[7983]<=26'd23451025;
ROM1[7984]<=26'd1971212; ROM2[7984]<=26'd11124348; ROM3[7984]<=26'd9722884; ROM4[7984]<=26'd23446840;
ROM1[7985]<=26'd1967727; ROM2[7985]<=26'd11126809; ROM3[7985]<=26'd9726423; ROM4[7985]<=26'd23448583;
ROM1[7986]<=26'd1969864; ROM2[7986]<=26'd11137502; ROM3[7986]<=26'd9735779; ROM4[7986]<=26'd23458918;
ROM1[7987]<=26'd1968649; ROM2[7987]<=26'd11138642; ROM3[7987]<=26'd9737727; ROM4[7987]<=26'd23459896;
ROM1[7988]<=26'd1968460; ROM2[7988]<=26'd11133867; ROM3[7988]<=26'd9730737; ROM4[7988]<=26'd23454000;
ROM1[7989]<=26'd1980480; ROM2[7989]<=26'd11135427; ROM3[7989]<=26'd9726982; ROM4[7989]<=26'd23453397;
ROM1[7990]<=26'd1992504; ROM2[7990]<=26'd11138682; ROM3[7990]<=26'd9726670; ROM4[7990]<=26'd23456590;
ROM1[7991]<=26'd1989794; ROM2[7991]<=26'd11138085; ROM3[7991]<=26'd9729765; ROM4[7991]<=26'd23458458;
ROM1[7992]<=26'd1980168; ROM2[7992]<=26'd11135952; ROM3[7992]<=26'd9731917; ROM4[7992]<=26'd23458012;
ROM1[7993]<=26'd1975265; ROM2[7993]<=26'd11136283; ROM3[7993]<=26'd9737001; ROM4[7993]<=26'd23459615;
ROM1[7994]<=26'd1974130; ROM2[7994]<=26'd11139600; ROM3[7994]<=26'd9743539; ROM4[7994]<=26'd23463051;
ROM1[7995]<=26'd1969447; ROM2[7995]<=26'd11139159; ROM3[7995]<=26'd9743566; ROM4[7995]<=26'd23461381;
ROM1[7996]<=26'd1971569; ROM2[7996]<=26'd11140062; ROM3[7996]<=26'd9743036; ROM4[7996]<=26'd23461962;
ROM1[7997]<=26'd1980691; ROM2[7997]<=26'd11141535; ROM3[7997]<=26'd9737490; ROM4[7997]<=26'd23462665;
ROM1[7998]<=26'd1993408; ROM2[7998]<=26'd11142417; ROM3[7998]<=26'd9732323; ROM4[7998]<=26'd23460327;
ROM1[7999]<=26'd1999309; ROM2[7999]<=26'd11147118; ROM3[7999]<=26'd9737313; ROM4[7999]<=26'd23464091;
ROM1[8000]<=26'd1993660; ROM2[8000]<=26'd11147044; ROM3[8000]<=26'd9740708; ROM4[8000]<=26'd23465388;
ROM1[8001]<=26'd1986692; ROM2[8001]<=26'd11143870; ROM3[8001]<=26'd9742660; ROM4[8001]<=26'd23463843;
ROM1[8002]<=26'd1984822; ROM2[8002]<=26'd11145623; ROM3[8002]<=26'd9747200; ROM4[8002]<=26'd23466264;
ROM1[8003]<=26'd1971944; ROM2[8003]<=26'd11137970; ROM3[8003]<=26'd9740798; ROM4[8003]<=26'd23460035;
ROM1[8004]<=26'd1966641; ROM2[8004]<=26'd11131601; ROM3[8004]<=26'd9732673; ROM4[8004]<=26'd23454759;
ROM1[8005]<=26'd1980066; ROM2[8005]<=26'd11136945; ROM3[8005]<=26'd9734367; ROM4[8005]<=26'd23458168;
ROM1[8006]<=26'd1990872; ROM2[8006]<=26'd11135656; ROM3[8006]<=26'd9727561; ROM4[8006]<=26'd23456236;
ROM1[8007]<=26'd1994484; ROM2[8007]<=26'd11133593; ROM3[8007]<=26'd9722803; ROM4[8007]<=26'd23454568;
ROM1[8008]<=26'd1993723; ROM2[8008]<=26'd11138801; ROM3[8008]<=26'd9729711; ROM4[8008]<=26'd23459474;
ROM1[8009]<=26'd1986670; ROM2[8009]<=26'd11140760; ROM3[8009]<=26'd9734412; ROM4[8009]<=26'd23461609;
ROM1[8010]<=26'd1982391; ROM2[8010]<=26'd11140790; ROM3[8010]<=26'd9738052; ROM4[8010]<=26'd23462464;
ROM1[8011]<=26'd1977819; ROM2[8011]<=26'd11140312; ROM3[8011]<=26'd9742515; ROM4[8011]<=26'd23464594;
ROM1[8012]<=26'd1977223; ROM2[8012]<=26'd11140640; ROM3[8012]<=26'd9744611; ROM4[8012]<=26'd23465363;
ROM1[8013]<=26'd1981693; ROM2[8013]<=26'd11141208; ROM3[8013]<=26'd9743570; ROM4[8013]<=26'd23465266;
ROM1[8014]<=26'd1991973; ROM2[8014]<=26'd11142609; ROM3[8014]<=26'd9740852; ROM4[8014]<=26'd23466104;
ROM1[8015]<=26'd2002406; ROM2[8015]<=26'd11145661; ROM3[8015]<=26'd9737019; ROM4[8015]<=26'd23466675;
ROM1[8016]<=26'd2001682; ROM2[8016]<=26'd11144824; ROM3[8016]<=26'd9737674; ROM4[8016]<=26'd23467114;
ROM1[8017]<=26'd1993595; ROM2[8017]<=26'd11143044; ROM3[8017]<=26'd9741106; ROM4[8017]<=26'd23468312;
ROM1[8018]<=26'd1985275; ROM2[8018]<=26'd11141645; ROM3[8018]<=26'd9744625; ROM4[8018]<=26'd23469259;
ROM1[8019]<=26'd1979852; ROM2[8019]<=26'd11139654; ROM3[8019]<=26'd9748691; ROM4[8019]<=26'd23469880;
ROM1[8020]<=26'd1976389; ROM2[8020]<=26'd11141247; ROM3[8020]<=26'd9752528; ROM4[8020]<=26'd23471883;
ROM1[8021]<=26'd1978674; ROM2[8021]<=26'd11142273; ROM3[8021]<=26'd9751214; ROM4[8021]<=26'd23472062;
ROM1[8022]<=26'd1988645; ROM2[8022]<=26'd11141378; ROM3[8022]<=26'd9747609; ROM4[8022]<=26'd23470293;
ROM1[8023]<=26'd2001996; ROM2[8023]<=26'd11143185; ROM3[8023]<=26'd9744653; ROM4[8023]<=26'd23471274;
ROM1[8024]<=26'd2003754; ROM2[8024]<=26'd11143625; ROM3[8024]<=26'd9745518; ROM4[8024]<=26'd23474504;
ROM1[8025]<=26'd2005103; ROM2[8025]<=26'd11151326; ROM3[8025]<=26'd9756108; ROM4[8025]<=26'd23481920;
ROM1[8026]<=26'd2000555; ROM2[8026]<=26'd11154493; ROM3[8026]<=26'd9761458; ROM4[8026]<=26'd23484980;
ROM1[8027]<=26'd1984778; ROM2[8027]<=26'd11144361; ROM3[8027]<=26'd9756226; ROM4[8027]<=26'd23477481;
ROM1[8028]<=26'd1976497; ROM2[8028]<=26'd11140561; ROM3[8028]<=26'd9755157; ROM4[8028]<=26'd23474510;
ROM1[8029]<=26'd1972727; ROM2[8029]<=26'd11134879; ROM3[8029]<=26'd9752344; ROM4[8029]<=26'd23471845;
ROM1[8030]<=26'd1978115; ROM2[8030]<=26'd11132365; ROM3[8030]<=26'd9747238; ROM4[8030]<=26'd23468933;
ROM1[8031]<=26'd1996052; ROM2[8031]<=26'd11139447; ROM3[8031]<=26'd9744751; ROM4[8031]<=26'd23472909;
ROM1[8032]<=26'd2003909; ROM2[8032]<=26'd11142886; ROM3[8032]<=26'd9746572; ROM4[8032]<=26'd23475451;
ROM1[8033]<=26'd2002527; ROM2[8033]<=26'd11146662; ROM3[8033]<=26'd9752906; ROM4[8033]<=26'd23480778;
ROM1[8034]<=26'd1994307; ROM2[8034]<=26'd11146983; ROM3[8034]<=26'd9755516; ROM4[8034]<=26'd23482101;
ROM1[8035]<=26'd1984510; ROM2[8035]<=26'd11142260; ROM3[8035]<=26'd9753178; ROM4[8035]<=26'd23476954;
ROM1[8036]<=26'd1975030; ROM2[8036]<=26'd11139299; ROM3[8036]<=26'd9750536; ROM4[8036]<=26'd23472009;
ROM1[8037]<=26'd1968450; ROM2[8037]<=26'd11135835; ROM3[8037]<=26'd9746022; ROM4[8037]<=26'd23465184;
ROM1[8038]<=26'd1980493; ROM2[8038]<=26'd11142855; ROM3[8038]<=26'd9747577; ROM4[8038]<=26'd23469588;
ROM1[8039]<=26'd1999563; ROM2[8039]<=26'd11150280; ROM3[8039]<=26'd9747372; ROM4[8039]<=26'd23475128;
ROM1[8040]<=26'd2003262; ROM2[8040]<=26'd11144137; ROM3[8040]<=26'd9736792; ROM4[8040]<=26'd23468931;
ROM1[8041]<=26'd1996802; ROM2[8041]<=26'd11139234; ROM3[8041]<=26'd9732006; ROM4[8041]<=26'd23463822;
ROM1[8042]<=26'd1984767; ROM2[8042]<=26'd11134503; ROM3[8042]<=26'd9731744; ROM4[8042]<=26'd23459160;
ROM1[8043]<=26'd1978576; ROM2[8043]<=26'd11134500; ROM3[8043]<=26'd9734383; ROM4[8043]<=26'd23459281;
ROM1[8044]<=26'd1977048; ROM2[8044]<=26'd11139430; ROM3[8044]<=26'd9739420; ROM4[8044]<=26'd23463733;
ROM1[8045]<=26'd1973629; ROM2[8045]<=26'd11141117; ROM3[8045]<=26'd9741743; ROM4[8045]<=26'd23464707;
ROM1[8046]<=26'd1978908; ROM2[8046]<=26'd11141526; ROM3[8046]<=26'd9741028; ROM4[8046]<=26'd23464940;
ROM1[8047]<=26'd1996041; ROM2[8047]<=26'd11147769; ROM3[8047]<=26'd9742585; ROM4[8047]<=26'd23469776;
ROM1[8048]<=26'd2010065; ROM2[8048]<=26'd11151883; ROM3[8048]<=26'd9740734; ROM4[8048]<=26'd23470730;
ROM1[8049]<=26'd2006034; ROM2[8049]<=26'd11147529; ROM3[8049]<=26'd9736185; ROM4[8049]<=26'd23466231;
ROM1[8050]<=26'd1994539; ROM2[8050]<=26'd11144639; ROM3[8050]<=26'd9735572; ROM4[8050]<=26'd23463133;
ROM1[8051]<=26'd1984644; ROM2[8051]<=26'd11142380; ROM3[8051]<=26'd9738130; ROM4[8051]<=26'd23461542;
ROM1[8052]<=26'd1978627; ROM2[8052]<=26'd11140946; ROM3[8052]<=26'd9742035; ROM4[8052]<=26'd23463013;
ROM1[8053]<=26'd1975398; ROM2[8053]<=26'd11143716; ROM3[8053]<=26'd9747898; ROM4[8053]<=26'd23466758;
ROM1[8054]<=26'd1979505; ROM2[8054]<=26'd11147991; ROM3[8054]<=26'd9751640; ROM4[8054]<=26'd23470790;
ROM1[8055]<=26'd1988026; ROM2[8055]<=26'd11148959; ROM3[8055]<=26'd9749849; ROM4[8055]<=26'd23470001;
ROM1[8056]<=26'd2003088; ROM2[8056]<=26'd11150864; ROM3[8056]<=26'd9748054; ROM4[8056]<=26'd23470506;
ROM1[8057]<=26'd2014252; ROM2[8057]<=26'd11155216; ROM3[8057]<=26'd9750141; ROM4[8057]<=26'd23476589;
ROM1[8058]<=26'd2004942; ROM2[8058]<=26'd11153079; ROM3[8058]<=26'd9750012; ROM4[8058]<=26'd23474245;
ROM1[8059]<=26'd1988418; ROM2[8059]<=26'd11144316; ROM3[8059]<=26'd9747168; ROM4[8059]<=26'd23468968;
ROM1[8060]<=26'd1980681; ROM2[8060]<=26'd11139944; ROM3[8060]<=26'd9746318; ROM4[8060]<=26'd23468121;
ROM1[8061]<=26'd1980435; ROM2[8061]<=26'd11143844; ROM3[8061]<=26'd9752858; ROM4[8061]<=26'd23472865;
ROM1[8062]<=26'd1994267; ROM2[8062]<=26'd11156214; ROM3[8062]<=26'd9767103; ROM4[8062]<=26'd23488324;
ROM1[8063]<=26'd2003114; ROM2[8063]<=26'd11161179; ROM3[8063]<=26'd9769831; ROM4[8063]<=26'd23492464;
ROM1[8064]<=26'd2010805; ROM2[8064]<=26'd11157643; ROM3[8064]<=26'd9760345; ROM4[8064]<=26'd23486462;
ROM1[8065]<=26'd2016766; ROM2[8065]<=26'd11154635; ROM3[8065]<=26'd9752389; ROM4[8065]<=26'd23483328;
ROM1[8066]<=26'd2008517; ROM2[8066]<=26'd11149745; ROM3[8066]<=26'd9748491; ROM4[8066]<=26'd23478816;
ROM1[8067]<=26'd2002522; ROM2[8067]<=26'd11150515; ROM3[8067]<=26'd9752414; ROM4[8067]<=26'd23480040;
ROM1[8068]<=26'd2001421; ROM2[8068]<=26'd11155625; ROM3[8068]<=26'd9763656; ROM4[8068]<=26'd23486879;
ROM1[8069]<=26'd1997790; ROM2[8069]<=26'd11156731; ROM3[8069]<=26'd9769525; ROM4[8069]<=26'd23489126;
ROM1[8070]<=26'd1991304; ROM2[8070]<=26'd11152167; ROM3[8070]<=26'd9769325; ROM4[8070]<=26'd23487345;
ROM1[8071]<=26'd1994215; ROM2[8071]<=26'd11152871; ROM3[8071]<=26'd9770797; ROM4[8071]<=26'd23488395;
ROM1[8072]<=26'd2005617; ROM2[8072]<=26'd11157392; ROM3[8072]<=26'd9768032; ROM4[8072]<=26'd23490281;
ROM1[8073]<=26'd2015842; ROM2[8073]<=26'd11155661; ROM3[8073]<=26'd9759891; ROM4[8073]<=26'd23488720;
ROM1[8074]<=26'd2015555; ROM2[8074]<=26'd11153239; ROM3[8074]<=26'd9756796; ROM4[8074]<=26'd23485683;
ROM1[8075]<=26'd2007765; ROM2[8075]<=26'd11150463; ROM3[8075]<=26'd9758430; ROM4[8075]<=26'd23484265;
ROM1[8076]<=26'd1999934; ROM2[8076]<=26'd11148353; ROM3[8076]<=26'd9760379; ROM4[8076]<=26'd23483914;
ROM1[8077]<=26'd1996925; ROM2[8077]<=26'd11150365; ROM3[8077]<=26'd9764678; ROM4[8077]<=26'd23486837;
ROM1[8078]<=26'd1998630; ROM2[8078]<=26'd11157113; ROM3[8078]<=26'd9772002; ROM4[8078]<=26'd23495220;
ROM1[8079]<=26'd2002117; ROM2[8079]<=26'd11160954; ROM3[8079]<=26'd9771748; ROM4[8079]<=26'd23497589;
ROM1[8080]<=26'd2000981; ROM2[8080]<=26'd11153524; ROM3[8080]<=26'd9760099; ROM4[8080]<=26'd23488629;
ROM1[8081]<=26'd2007802; ROM2[8081]<=26'd11150689; ROM3[8081]<=26'd9750909; ROM4[8081]<=26'd23483956;
ROM1[8082]<=26'd2009681; ROM2[8082]<=26'd11148894; ROM3[8082]<=26'd9746090; ROM4[8082]<=26'd23480970;
ROM1[8083]<=26'd2005584; ROM2[8083]<=26'd11148435; ROM3[8083]<=26'd9747027; ROM4[8083]<=26'd23482712;
ROM1[8084]<=26'd2006075; ROM2[8084]<=26'd11154699; ROM3[8084]<=26'd9757681; ROM4[8084]<=26'd23490590;
ROM1[8085]<=26'd2006088; ROM2[8085]<=26'd11158213; ROM3[8085]<=26'd9766381; ROM4[8085]<=26'd23494750;
ROM1[8086]<=26'd1993291; ROM2[8086]<=26'd11152799; ROM3[8086]<=26'd9763934; ROM4[8086]<=26'd23489992;
ROM1[8087]<=26'd1974191; ROM2[8087]<=26'd11139004; ROM3[8087]<=26'd9749082; ROM4[8087]<=26'd23473787;
ROM1[8088]<=26'd1977781; ROM2[8088]<=26'd11138085; ROM3[8088]<=26'd9741885; ROM4[8088]<=26'd23467829;
ROM1[8089]<=26'd1992601; ROM2[8089]<=26'd11143484; ROM3[8089]<=26'd9738149; ROM4[8089]<=26'd23470137;
ROM1[8090]<=26'd1998957; ROM2[8090]<=26'd11140484; ROM3[8090]<=26'd9731301; ROM4[8090]<=26'd23466448;
ROM1[8091]<=26'd2000085; ROM2[8091]<=26'd11143318; ROM3[8091]<=26'd9735736; ROM4[8091]<=26'd23469106;
ROM1[8092]<=26'd1991833; ROM2[8092]<=26'd11142778; ROM3[8092]<=26'd9739880; ROM4[8092]<=26'd23471336;
ROM1[8093]<=26'd1976502; ROM2[8093]<=26'd11134852; ROM3[8093]<=26'd9737165; ROM4[8093]<=26'd23464817;
ROM1[8094]<=26'd1970196; ROM2[8094]<=26'd11133040; ROM3[8094]<=26'd9739343; ROM4[8094]<=26'd23463394;
ROM1[8095]<=26'd1969584; ROM2[8095]<=26'd11134589; ROM3[8095]<=26'd9743509; ROM4[8095]<=26'd23465219;
ROM1[8096]<=26'd1975492; ROM2[8096]<=26'd11140914; ROM3[8096]<=26'd9746824; ROM4[8096]<=26'd23470072;
ROM1[8097]<=26'd1985649; ROM2[8097]<=26'd11142107; ROM3[8097]<=26'd9741889; ROM4[8097]<=26'd23468252;
ROM1[8098]<=26'd1996041; ROM2[8098]<=26'd11141625; ROM3[8098]<=26'd9734139; ROM4[8098]<=26'd23465180;
ROM1[8099]<=26'd1994824; ROM2[8099]<=26'd11140637; ROM3[8099]<=26'd9731111; ROM4[8099]<=26'd23464488;
ROM1[8100]<=26'd1983128; ROM2[8100]<=26'd11134425; ROM3[8100]<=26'd9728472; ROM4[8100]<=26'd23458520;
ROM1[8101]<=26'd1976008; ROM2[8101]<=26'd11133292; ROM3[8101]<=26'd9732331; ROM4[8101]<=26'd23458563;
ROM1[8102]<=26'd1973926; ROM2[8102]<=26'd11135636; ROM3[8102]<=26'd9736235; ROM4[8102]<=26'd23462120;
ROM1[8103]<=26'd1969577; ROM2[8103]<=26'd11137189; ROM3[8103]<=26'd9739826; ROM4[8103]<=26'd23463790;
ROM1[8104]<=26'd1970436; ROM2[8104]<=26'd11138191; ROM3[8104]<=26'd9740402; ROM4[8104]<=26'd23464265;
ROM1[8105]<=26'd1980923; ROM2[8105]<=26'd11141716; ROM3[8105]<=26'd9740330; ROM4[8105]<=26'd23465744;
ROM1[8106]<=26'd1994450; ROM2[8106]<=26'd11143560; ROM3[8106]<=26'd9735805; ROM4[8106]<=26'd23466036;
ROM1[8107]<=26'd1998554; ROM2[8107]<=26'd11143107; ROM3[8107]<=26'd9733458; ROM4[8107]<=26'd23466397;
ROM1[8108]<=26'd1994171; ROM2[8108]<=26'd11143264; ROM3[8108]<=26'd9735407; ROM4[8108]<=26'd23467570;
ROM1[8109]<=26'd1986033; ROM2[8109]<=26'd11141826; ROM3[8109]<=26'd9736896; ROM4[8109]<=26'd23467819;
ROM1[8110]<=26'd1978094; ROM2[8110]<=26'd11140556; ROM3[8110]<=26'd9740051; ROM4[8110]<=26'd23466698;
ROM1[8111]<=26'd1973129; ROM2[8111]<=26'd11140931; ROM3[8111]<=26'd9744266; ROM4[8111]<=26'd23468032;
ROM1[8112]<=26'd1970917; ROM2[8112]<=26'd11139985; ROM3[8112]<=26'd9744658; ROM4[8112]<=26'd23467911;
ROM1[8113]<=26'd1975070; ROM2[8113]<=26'd11138612; ROM3[8113]<=26'd9741918; ROM4[8113]<=26'd23465749;
ROM1[8114]<=26'd1991264; ROM2[8114]<=26'd11144366; ROM3[8114]<=26'd9742402; ROM4[8114]<=26'd23468341;
ROM1[8115]<=26'd2000377; ROM2[8115]<=26'd11147585; ROM3[8115]<=26'd9740324; ROM4[8115]<=26'd23468351;
ROM1[8116]<=26'd1994667; ROM2[8116]<=26'd11146187; ROM3[8116]<=26'd9738841; ROM4[8116]<=26'd23465224;
ROM1[8117]<=26'd1986241; ROM2[8117]<=26'd11145011; ROM3[8117]<=26'd9740983; ROM4[8117]<=26'd23464233;
ROM1[8118]<=26'd1977742; ROM2[8118]<=26'd11141802; ROM3[8118]<=26'd9742052; ROM4[8118]<=26'd23463914;
ROM1[8119]<=26'd1971659; ROM2[8119]<=26'd11140268; ROM3[8119]<=26'd9742747; ROM4[8119]<=26'd23463897;
ROM1[8120]<=26'd1967531; ROM2[8120]<=26'd11141272; ROM3[8120]<=26'd9746437; ROM4[8120]<=26'd23465875;
ROM1[8121]<=26'd1970309; ROM2[8121]<=26'd11142649; ROM3[8121]<=26'd9746385; ROM4[8121]<=26'd23466607;
ROM1[8122]<=26'd1981613; ROM2[8122]<=26'd11145748; ROM3[8122]<=26'd9742214; ROM4[8122]<=26'd23467445;
ROM1[8123]<=26'd1997640; ROM2[8123]<=26'd11150029; ROM3[8123]<=26'd9740989; ROM4[8123]<=26'd23472242;
ROM1[8124]<=26'd2001966; ROM2[8124]<=26'd11151353; ROM3[8124]<=26'd9743782; ROM4[8124]<=26'd23475111;
ROM1[8125]<=26'd1998013; ROM2[8125]<=26'd11152016; ROM3[8125]<=26'd9749143; ROM4[8125]<=26'd23478976;
ROM1[8126]<=26'd1992839; ROM2[8126]<=26'd11152436; ROM3[8126]<=26'd9755554; ROM4[8126]<=26'd23481931;
ROM1[8127]<=26'd1984055; ROM2[8127]<=26'd11147622; ROM3[8127]<=26'd9755636; ROM4[8127]<=26'd23478460;
ROM1[8128]<=26'd1973357; ROM2[8128]<=26'd11139756; ROM3[8128]<=26'd9752388; ROM4[8128]<=26'd23474637;
ROM1[8129]<=26'd1972160; ROM2[8129]<=26'd11137044; ROM3[8129]<=26'd9750258; ROM4[8129]<=26'd23472808;
ROM1[8130]<=26'd1978301; ROM2[8130]<=26'd11135573; ROM3[8130]<=26'd9746692; ROM4[8130]<=26'd23470955;
ROM1[8131]<=26'd1992786; ROM2[8131]<=26'd11137674; ROM3[8131]<=26'd9742389; ROM4[8131]<=26'd23473182;
ROM1[8132]<=26'd2000221; ROM2[8132]<=26'd11139467; ROM3[8132]<=26'd9742607; ROM4[8132]<=26'd23475682;
ROM1[8133]<=26'd1992338; ROM2[8133]<=26'd11136211; ROM3[8133]<=26'd9741673; ROM4[8133]<=26'd23471629;
ROM1[8134]<=26'd1984451; ROM2[8134]<=26'd11133371; ROM3[8134]<=26'd9744774; ROM4[8134]<=26'd23468720;
ROM1[8135]<=26'd1982725; ROM2[8135]<=26'd11135715; ROM3[8135]<=26'd9750559; ROM4[8135]<=26'd23470925;
ROM1[8136]<=26'd1982853; ROM2[8136]<=26'd11144305; ROM3[8136]<=26'd9756820; ROM4[8136]<=26'd23476439;
ROM1[8137]<=26'd1976672; ROM2[8137]<=26'd11140473; ROM3[8137]<=26'd9753466; ROM4[8137]<=26'd23471923;
ROM1[8138]<=26'd1974375; ROM2[8138]<=26'd11132233; ROM3[8138]<=26'd9742910; ROM4[8138]<=26'd23464091;
ROM1[8139]<=26'd1987552; ROM2[8139]<=26'd11135810; ROM3[8139]<=26'd9738337; ROM4[8139]<=26'd23463882;
ROM1[8140]<=26'd1990933; ROM2[8140]<=26'd11132187; ROM3[8140]<=26'd9729957; ROM4[8140]<=26'd23458106;
ROM1[8141]<=26'd1986401; ROM2[8141]<=26'd11131334; ROM3[8141]<=26'd9729339; ROM4[8141]<=26'd23458811;
ROM1[8142]<=26'd1984318; ROM2[8142]<=26'd11137749; ROM3[8142]<=26'd9735727; ROM4[8142]<=26'd23465175;
ROM1[8143]<=26'd1977581; ROM2[8143]<=26'd11138676; ROM3[8143]<=26'd9741159; ROM4[8143]<=26'd23466387;
ROM1[8144]<=26'd1973917; ROM2[8144]<=26'd11137971; ROM3[8144]<=26'd9746084; ROM4[8144]<=26'd23469318;
ROM1[8145]<=26'd1969753; ROM2[8145]<=26'd11138150; ROM3[8145]<=26'd9747712; ROM4[8145]<=26'd23469793;
ROM1[8146]<=26'd1969677; ROM2[8146]<=26'd11137704; ROM3[8146]<=26'd9745432; ROM4[8146]<=26'd23468718;
ROM1[8147]<=26'd1975947; ROM2[8147]<=26'd11135486; ROM3[8147]<=26'd9737837; ROM4[8147]<=26'd23465588;
ROM1[8148]<=26'd1984612; ROM2[8148]<=26'd11133954; ROM3[8148]<=26'd9730025; ROM4[8148]<=26'd23461821;
ROM1[8149]<=26'd1987009; ROM2[8149]<=26'd11134842; ROM3[8149]<=26'd9729475; ROM4[8149]<=26'd23462298;
ROM1[8150]<=26'd1981742; ROM2[8150]<=26'd11135871; ROM3[8150]<=26'd9732266; ROM4[8150]<=26'd23464192;
ROM1[8151]<=26'd1975600; ROM2[8151]<=26'd11136160; ROM3[8151]<=26'd9736914; ROM4[8151]<=26'd23464745;
ROM1[8152]<=26'd1976653; ROM2[8152]<=26'd11141978; ROM3[8152]<=26'd9746126; ROM4[8152]<=26'd23469971;
ROM1[8153]<=26'd1976777; ROM2[8153]<=26'd11148476; ROM3[8153]<=26'd9753439; ROM4[8153]<=26'd23475392;
ROM1[8154]<=26'd1972790; ROM2[8154]<=26'd11144810; ROM3[8154]<=26'd9748619; ROM4[8154]<=26'd23469578;
ROM1[8155]<=26'd1973325; ROM2[8155]<=26'd11137361; ROM3[8155]<=26'd9737210; ROM4[8155]<=26'd23460879;
ROM1[8156]<=26'd1984154; ROM2[8156]<=26'd11135470; ROM3[8156]<=26'd9728420; ROM4[8156]<=26'd23456824;
ROM1[8157]<=26'd1987368; ROM2[8157]<=26'd11133620; ROM3[8157]<=26'd9721568; ROM4[8157]<=26'd23454505;
ROM1[8158]<=26'd1980291; ROM2[8158]<=26'd11131214; ROM3[8158]<=26'd9721572; ROM4[8158]<=26'd23453976;
ROM1[8159]<=26'd1973755; ROM2[8159]<=26'd11130762; ROM3[8159]<=26'd9727844; ROM4[8159]<=26'd23455406;
ROM1[8160]<=26'd1965786; ROM2[8160]<=26'd11128182; ROM3[8160]<=26'd9726956; ROM4[8160]<=26'd23453679;
ROM1[8161]<=26'd1958636; ROM2[8161]<=26'd11126187; ROM3[8161]<=26'd9729738; ROM4[8161]<=26'd23452610;
ROM1[8162]<=26'd1963723; ROM2[8162]<=26'd11133364; ROM3[8162]<=26'd9737567; ROM4[8162]<=26'd23459173;
ROM1[8163]<=26'd1975664; ROM2[8163]<=26'd11140392; ROM3[8163]<=26'd9739707; ROM4[8163]<=26'd23464677;
ROM1[8164]<=26'd1986978; ROM2[8164]<=26'd11139515; ROM3[8164]<=26'd9734431; ROM4[8164]<=26'd23462541;
ROM1[8165]<=26'd1994486; ROM2[8165]<=26'd11138748; ROM3[8165]<=26'd9728827; ROM4[8165]<=26'd23459869;
ROM1[8166]<=26'd1984572; ROM2[8166]<=26'd11132001; ROM3[8166]<=26'd9721259; ROM4[8166]<=26'd23451802;
ROM1[8167]<=26'd1972987; ROM2[8167]<=26'd11125444; ROM3[8167]<=26'd9718215; ROM4[8167]<=26'd23445243;
ROM1[8168]<=26'd1964245; ROM2[8168]<=26'd11123798; ROM3[8168]<=26'd9721052; ROM4[8168]<=26'd23443109;
ROM1[8169]<=26'd1957858; ROM2[8169]<=26'd11122027; ROM3[8169]<=26'd9721117; ROM4[8169]<=26'd23440859;
ROM1[8170]<=26'd1956738; ROM2[8170]<=26'd11122126; ROM3[8170]<=26'd9723027; ROM4[8170]<=26'd23440701;
ROM1[8171]<=26'd1957584; ROM2[8171]<=26'd11122670; ROM3[8171]<=26'd9720200; ROM4[8171]<=26'd23440168;
ROM1[8172]<=26'd1968069; ROM2[8172]<=26'd11124346; ROM3[8172]<=26'd9714334; ROM4[8172]<=26'd23440216;
ROM1[8173]<=26'd1981578; ROM2[8173]<=26'd11127788; ROM3[8173]<=26'd9712389; ROM4[8173]<=26'd23443283;
ROM1[8174]<=26'd1982158; ROM2[8174]<=26'd11128304; ROM3[8174]<=26'd9714423; ROM4[8174]<=26'd23445175;
ROM1[8175]<=26'd1976804; ROM2[8175]<=26'd11127538; ROM3[8175]<=26'd9716143; ROM4[8175]<=26'd23446299;
ROM1[8176]<=26'd1972608; ROM2[8176]<=26'd11129733; ROM3[8176]<=26'd9721145; ROM4[8176]<=26'd23449209;
ROM1[8177]<=26'd1968005; ROM2[8177]<=26'd11131834; ROM3[8177]<=26'd9725826; ROM4[8177]<=26'd23451637;
ROM1[8178]<=26'd1966213; ROM2[8178]<=26'd11135558; ROM3[8178]<=26'd9731189; ROM4[8178]<=26'd23456968;
ROM1[8179]<=26'd1972272; ROM2[8179]<=26'd11141998; ROM3[8179]<=26'd9740745; ROM4[8179]<=26'd23463245;
ROM1[8180]<=26'd1984220; ROM2[8180]<=26'd11146155; ROM3[8180]<=26'd9743014; ROM4[8180]<=26'd23467124;
ROM1[8181]<=26'd2000568; ROM2[8181]<=26'd11148213; ROM3[8181]<=26'd9739352; ROM4[8181]<=26'd23470560;
ROM1[8182]<=26'd2003757; ROM2[8182]<=26'd11146233; ROM3[8182]<=26'd9738161; ROM4[8182]<=26'd23469788;
ROM1[8183]<=26'd1998221; ROM2[8183]<=26'd11143792; ROM3[8183]<=26'd9741371; ROM4[8183]<=26'd23471087;
ROM1[8184]<=26'd1992887; ROM2[8184]<=26'd11145779; ROM3[8184]<=26'd9748016; ROM4[8184]<=26'd23475603;
ROM1[8185]<=26'd1984899; ROM2[8185]<=26'd11140488; ROM3[8185]<=26'd9748922; ROM4[8185]<=26'd23470979;
ROM1[8186]<=26'd1978928; ROM2[8186]<=26'd11139312; ROM3[8186]<=26'd9751675; ROM4[8186]<=26'd23472259;
ROM1[8187]<=26'd1974405; ROM2[8187]<=26'd11137575; ROM3[8187]<=26'd9751468; ROM4[8187]<=26'd23471061;
ROM1[8188]<=26'd1980226; ROM2[8188]<=26'd11134579; ROM3[8188]<=26'd9748841; ROM4[8188]<=26'd23469285;
ROM1[8189]<=26'd1996574; ROM2[8189]<=26'd11138971; ROM3[8189]<=26'd9748079; ROM4[8189]<=26'd23474193;
ROM1[8190]<=26'd2005840; ROM2[8190]<=26'd11139162; ROM3[8190]<=26'd9744264; ROM4[8190]<=26'd23471666;
ROM1[8191]<=26'd2005428; ROM2[8191]<=26'd11139445; ROM3[8191]<=26'd9744205; ROM4[8191]<=26'd23471378;
ROM1[8192]<=26'd1994537; ROM2[8192]<=26'd11136411; ROM3[8192]<=26'd9744574; ROM4[8192]<=26'd23469929;
ROM1[8193]<=26'd1987286; ROM2[8193]<=26'd11137068; ROM3[8193]<=26'd9749538; ROM4[8193]<=26'd23472061;
ROM1[8194]<=26'd1986152; ROM2[8194]<=26'd11141335; ROM3[8194]<=26'd9754295; ROM4[8194]<=26'd23476788;
ROM1[8195]<=26'd1977003; ROM2[8195]<=26'd11135605; ROM3[8195]<=26'd9750025; ROM4[8195]<=26'd23469968;
ROM1[8196]<=26'd1975706; ROM2[8196]<=26'd11131353; ROM3[8196]<=26'd9744074; ROM4[8196]<=26'd23464101;
ROM1[8197]<=26'd1985136; ROM2[8197]<=26'd11131696; ROM3[8197]<=26'd9736683; ROM4[8197]<=26'd23461555;
ROM1[8198]<=26'd1995296; ROM2[8198]<=26'd11129347; ROM3[8198]<=26'd9729368; ROM4[8198]<=26'd23458544;
ROM1[8199]<=26'd1996868; ROM2[8199]<=26'd11131859; ROM3[8199]<=26'd9731248; ROM4[8199]<=26'd23460613;
ROM1[8200]<=26'd1991050; ROM2[8200]<=26'd11132738; ROM3[8200]<=26'd9734803; ROM4[8200]<=26'd23460335;
ROM1[8201]<=26'd1985189; ROM2[8201]<=26'd11132324; ROM3[8201]<=26'd9741066; ROM4[8201]<=26'd23462533;
ROM1[8202]<=26'd1985920; ROM2[8202]<=26'd11139314; ROM3[8202]<=26'd9751296; ROM4[8202]<=26'd23470278;
ROM1[8203]<=26'd1981403; ROM2[8203]<=26'd11140352; ROM3[8203]<=26'd9753004; ROM4[8203]<=26'd23471735;
ROM1[8204]<=26'd1974995; ROM2[8204]<=26'd11135453; ROM3[8204]<=26'd9748386; ROM4[8204]<=26'd23467614;
ROM1[8205]<=26'd1983023; ROM2[8205]<=26'd11137828; ROM3[8205]<=26'd9746993; ROM4[8205]<=26'd23467584;
ROM1[8206]<=26'd1997870; ROM2[8206]<=26'd11140283; ROM3[8206]<=26'd9742375; ROM4[8206]<=26'd23468104;
ROM1[8207]<=26'd1999758; ROM2[8207]<=26'd11137877; ROM3[8207]<=26'd9735222; ROM4[8207]<=26'd23466888;
ROM1[8208]<=26'd1993272; ROM2[8208]<=26'd11137933; ROM3[8208]<=26'd9736690; ROM4[8208]<=26'd23468152;
ROM1[8209]<=26'd1981195; ROM2[8209]<=26'd11133683; ROM3[8209]<=26'd9735673; ROM4[8209]<=26'd23464485;
ROM1[8210]<=26'd1970496; ROM2[8210]<=26'd11129235; ROM3[8210]<=26'd9734276; ROM4[8210]<=26'd23459670;
ROM1[8211]<=26'd1969499; ROM2[8211]<=26'd11133527; ROM3[8211]<=26'd9741850; ROM4[8211]<=26'd23463268;
ROM1[8212]<=26'd1975133; ROM2[8212]<=26'd11139835; ROM3[8212]<=26'd9746237; ROM4[8212]<=26'd23468675;
ROM1[8213]<=26'd1981371; ROM2[8213]<=26'd11140669; ROM3[8213]<=26'd9741988; ROM4[8213]<=26'd23467149;
ROM1[8214]<=26'd1988270; ROM2[8214]<=26'd11137492; ROM3[8214]<=26'd9733858; ROM4[8214]<=26'd23462768;
ROM1[8215]<=26'd1993335; ROM2[8215]<=26'd11136165; ROM3[8215]<=26'd9730129; ROM4[8215]<=26'd23460209;
ROM1[8216]<=26'd1994357; ROM2[8216]<=26'd11139278; ROM3[8216]<=26'd9737186; ROM4[8216]<=26'd23465453;
ROM1[8217]<=26'd1988186; ROM2[8217]<=26'd11139673; ROM3[8217]<=26'd9743404; ROM4[8217]<=26'd23469037;
ROM1[8218]<=26'd1973108; ROM2[8218]<=26'd11129403; ROM3[8218]<=26'd9737627; ROM4[8218]<=26'd23461635;
ROM1[8219]<=26'd1969223; ROM2[8219]<=26'd11127341; ROM3[8219]<=26'd9739974; ROM4[8219]<=26'd23462694;
ROM1[8220]<=26'd1970534; ROM2[8220]<=26'd11130731; ROM3[8220]<=26'd9743983; ROM4[8220]<=26'd23467062;
ROM1[8221]<=26'd1971716; ROM2[8221]<=26'd11127371; ROM3[8221]<=26'd9742804; ROM4[8221]<=26'd23465923;
ROM1[8222]<=26'd1982346; ROM2[8222]<=26'd11129208; ROM3[8222]<=26'd9741934; ROM4[8222]<=26'd23465760;
ROM1[8223]<=26'd1993184; ROM2[8223]<=26'd11131247; ROM3[8223]<=26'd9735842; ROM4[8223]<=26'd23464821;
ROM1[8224]<=26'd1988926; ROM2[8224]<=26'd11125721; ROM3[8224]<=26'd9732189; ROM4[8224]<=26'd23460664;
ROM1[8225]<=26'd1982971; ROM2[8225]<=26'd11125067; ROM3[8225]<=26'd9733698; ROM4[8225]<=26'd23459899;
ROM1[8226]<=26'd1981874; ROM2[8226]<=26'd11131127; ROM3[8226]<=26'd9740122; ROM4[8226]<=26'd23465875;
ROM1[8227]<=26'd1976535; ROM2[8227]<=26'd11130271; ROM3[8227]<=26'd9742943; ROM4[8227]<=26'd23466784;
ROM1[8228]<=26'd1968841; ROM2[8228]<=26'd11129030; ROM3[8228]<=26'd9743647; ROM4[8228]<=26'd23465475;
ROM1[8229]<=26'd1969687; ROM2[8229]<=26'd11130044; ROM3[8229]<=26'd9743864; ROM4[8229]<=26'd23464886;
ROM1[8230]<=26'd1979906; ROM2[8230]<=26'd11130221; ROM3[8230]<=26'd9741613; ROM4[8230]<=26'd23464445;
ROM1[8231]<=26'd1994565; ROM2[8231]<=26'd11132139; ROM3[8231]<=26'd9736761; ROM4[8231]<=26'd23465672;
ROM1[8232]<=26'd1997740; ROM2[8232]<=26'd11131766; ROM3[8232]<=26'd9733630; ROM4[8232]<=26'd23464608;
ROM1[8233]<=26'd1991464; ROM2[8233]<=26'd11132343; ROM3[8233]<=26'd9734538; ROM4[8233]<=26'd23463686;
ROM1[8234]<=26'd1987293; ROM2[8234]<=26'd11135437; ROM3[8234]<=26'd9739552; ROM4[8234]<=26'd23467570;
ROM1[8235]<=26'd1980902; ROM2[8235]<=26'd11133776; ROM3[8235]<=26'd9742093; ROM4[8235]<=26'd23466331;
ROM1[8236]<=26'd1972584; ROM2[8236]<=26'd11129709; ROM3[8236]<=26'd9739334; ROM4[8236]<=26'd23461202;
ROM1[8237]<=26'd1969191; ROM2[8237]<=26'd11127586; ROM3[8237]<=26'd9737105; ROM4[8237]<=26'd23457760;
ROM1[8238]<=26'd1972208; ROM2[8238]<=26'd11127977; ROM3[8238]<=26'd9734436; ROM4[8238]<=26'd23455081;
ROM1[8239]<=26'd1985121; ROM2[8239]<=26'd11131380; ROM3[8239]<=26'd9729459; ROM4[8239]<=26'd23455496;
ROM1[8240]<=26'd1998822; ROM2[8240]<=26'd11137482; ROM3[8240]<=26'd9731265; ROM4[8240]<=26'd23459453;
ROM1[8241]<=26'd1998889; ROM2[8241]<=26'd11140128; ROM3[8241]<=26'd9735672; ROM4[8241]<=26'd23461899;
ROM1[8242]<=26'd1986491; ROM2[8242]<=26'd11134611; ROM3[8242]<=26'd9733854; ROM4[8242]<=26'd23457930;
ROM1[8243]<=26'd1974404; ROM2[8243]<=26'd11128636; ROM3[8243]<=26'd9732873; ROM4[8243]<=26'd23453397;
ROM1[8244]<=26'd1968614; ROM2[8244]<=26'd11129659; ROM3[8244]<=26'd9736867; ROM4[8244]<=26'd23454768;
ROM1[8245]<=26'd1968048; ROM2[8245]<=26'd11134217; ROM3[8245]<=26'd9745661; ROM4[8245]<=26'd23461883;
ROM1[8246]<=26'd1969106; ROM2[8246]<=26'd11132390; ROM3[8246]<=26'd9746412; ROM4[8246]<=26'd23462543;
ROM1[8247]<=26'd1979711; ROM2[8247]<=26'd11130751; ROM3[8247]<=26'd9742556; ROM4[8247]<=26'd23461018;
ROM1[8248]<=26'd1994538; ROM2[8248]<=26'd11131985; ROM3[8248]<=26'd9741535; ROM4[8248]<=26'd23463354;
ROM1[8249]<=26'd1986628; ROM2[8249]<=26'd11123862; ROM3[8249]<=26'd9733021; ROM4[8249]<=26'd23456988;
ROM1[8250]<=26'd1981410; ROM2[8250]<=26'd11123691; ROM3[8250]<=26'd9735594; ROM4[8250]<=26'd23457599;
ROM1[8251]<=26'd1980751; ROM2[8251]<=26'd11132060; ROM3[8251]<=26'd9747078; ROM4[8251]<=26'd23466019;
ROM1[8252]<=26'd1969527; ROM2[8252]<=26'd11128356; ROM3[8252]<=26'd9743734; ROM4[8252]<=26'd23462769;
ROM1[8253]<=26'd1961206; ROM2[8253]<=26'd11125235; ROM3[8253]<=26'd9741048; ROM4[8253]<=26'd23458568;
ROM1[8254]<=26'd1965035; ROM2[8254]<=26'd11127956; ROM3[8254]<=26'd9742833; ROM4[8254]<=26'd23462040;
ROM1[8255]<=26'd1976818; ROM2[8255]<=26'd11131835; ROM3[8255]<=26'd9741505; ROM4[8255]<=26'd23465592;
ROM1[8256]<=26'd1996683; ROM2[8256]<=26'd11139538; ROM3[8256]<=26'd9741739; ROM4[8256]<=26'd23471206;
ROM1[8257]<=26'd1999257; ROM2[8257]<=26'd11138141; ROM3[8257]<=26'd9737351; ROM4[8257]<=26'd23469648;
ROM1[8258]<=26'd1988155; ROM2[8258]<=26'd11132400; ROM3[8258]<=26'd9731967; ROM4[8258]<=26'd23462949;
ROM1[8259]<=26'd1981573; ROM2[8259]<=26'd11131817; ROM3[8259]<=26'd9735071; ROM4[8259]<=26'd23463929;
ROM1[8260]<=26'd1975832; ROM2[8260]<=26'd11129689; ROM3[8260]<=26'd9737049; ROM4[8260]<=26'd23464701;
ROM1[8261]<=26'd1972167; ROM2[8261]<=26'd11131130; ROM3[8261]<=26'd9742148; ROM4[8261]<=26'd23466365;
ROM1[8262]<=26'd1970081; ROM2[8262]<=26'd11130229; ROM3[8262]<=26'd9742598; ROM4[8262]<=26'd23465299;
ROM1[8263]<=26'd1971439; ROM2[8263]<=26'd11125341; ROM3[8263]<=26'd9736601; ROM4[8263]<=26'd23460909;
ROM1[8264]<=26'd1979822; ROM2[8264]<=26'd11124316; ROM3[8264]<=26'd9729331; ROM4[8264]<=26'd23456064;
ROM1[8265]<=26'd1995525; ROM2[8265]<=26'd11132272; ROM3[8265]<=26'd9730619; ROM4[8265]<=26'd23462934;
ROM1[8266]<=26'd2010212; ROM2[8266]<=26'd11149748; ROM3[8266]<=26'd9749407; ROM4[8266]<=26'd23482642;
ROM1[8267]<=26'd1999283; ROM2[8267]<=26'd11143864; ROM3[8267]<=26'd9750468; ROM4[8267]<=26'd23479996;
ROM1[8268]<=26'd1981881; ROM2[8268]<=26'd11130934; ROM3[8268]<=26'd9742779; ROM4[8268]<=26'd23468888;
ROM1[8269]<=26'd1975653; ROM2[8269]<=26'd11130158; ROM3[8269]<=26'd9745399; ROM4[8269]<=26'd23470013;
ROM1[8270]<=26'd1968270; ROM2[8270]<=26'd11127094; ROM3[8270]<=26'd9743452; ROM4[8270]<=26'd23467157;
ROM1[8271]<=26'd1972415; ROM2[8271]<=26'd11130479; ROM3[8271]<=26'd9742916; ROM4[8271]<=26'd23467879;
ROM1[8272]<=26'd1988337; ROM2[8272]<=26'd11137559; ROM3[8272]<=26'd9743944; ROM4[8272]<=26'd23473842;
ROM1[8273]<=26'd2000233; ROM2[8273]<=26'd11140640; ROM3[8273]<=26'd9741421; ROM4[8273]<=26'd23474943;
ROM1[8274]<=26'd1996589; ROM2[8274]<=26'd11136840; ROM3[8274]<=26'd9738014; ROM4[8274]<=26'd23471576;
ROM1[8275]<=26'd1989516; ROM2[8275]<=26'd11133991; ROM3[8275]<=26'd9738293; ROM4[8275]<=26'd23469878;
ROM1[8276]<=26'd1982460; ROM2[8276]<=26'd11133082; ROM3[8276]<=26'd9742012; ROM4[8276]<=26'd23470136;
ROM1[8277]<=26'd1975467; ROM2[8277]<=26'd11129250; ROM3[8277]<=26'd9742345; ROM4[8277]<=26'd23469041;
ROM1[8278]<=26'd1969865; ROM2[8278]<=26'd11129397; ROM3[8278]<=26'd9742966; ROM4[8278]<=26'd23469346;
ROM1[8279]<=26'd1972231; ROM2[8279]<=26'd11134144; ROM3[8279]<=26'd9744783; ROM4[8279]<=26'd23471149;
ROM1[8280]<=26'd1982097; ROM2[8280]<=26'd11136343; ROM3[8280]<=26'd9742234; ROM4[8280]<=26'd23471641;
ROM1[8281]<=26'd1995468; ROM2[8281]<=26'd11136951; ROM3[8281]<=26'd9736032; ROM4[8281]<=26'd23469955;
ROM1[8282]<=26'd1994597; ROM2[8282]<=26'd11132611; ROM3[8282]<=26'd9728822; ROM4[8282]<=26'd23464995;
ROM1[8283]<=26'd1986486; ROM2[8283]<=26'd11130324; ROM3[8283]<=26'd9727492; ROM4[8283]<=26'd23461418;
ROM1[8284]<=26'd1980148; ROM2[8284]<=26'd11130052; ROM3[8284]<=26'd9730629; ROM4[8284]<=26'd23460661;
ROM1[8285]<=26'd1974057; ROM2[8285]<=26'd11129212; ROM3[8285]<=26'd9732263; ROM4[8285]<=26'd23461277;
ROM1[8286]<=26'd1972273; ROM2[8286]<=26'd11132195; ROM3[8286]<=26'd9737171; ROM4[8286]<=26'd23464709;
ROM1[8287]<=26'd1971415; ROM2[8287]<=26'd11132436; ROM3[8287]<=26'd9740176; ROM4[8287]<=26'd23466521;
ROM1[8288]<=26'd1974851; ROM2[8288]<=26'd11132327; ROM3[8288]<=26'd9737793; ROM4[8288]<=26'd23468084;
ROM1[8289]<=26'd1989192; ROM2[8289]<=26'd11134070; ROM3[8289]<=26'd9734615; ROM4[8289]<=26'd23468421;
ROM1[8290]<=26'd2001121; ROM2[8290]<=26'd11137869; ROM3[8290]<=26'd9736042; ROM4[8290]<=26'd23469907;
ROM1[8291]<=26'd1998862; ROM2[8291]<=26'd11138843; ROM3[8291]<=26'd9738854; ROM4[8291]<=26'd23472108;
ROM1[8292]<=26'd1994255; ROM2[8292]<=26'd11141065; ROM3[8292]<=26'd9744586; ROM4[8292]<=26'd23474918;
ROM1[8293]<=26'd1991377; ROM2[8293]<=26'd11143210; ROM3[8293]<=26'd9750091; ROM4[8293]<=26'd23478151;
ROM1[8294]<=26'd1983111; ROM2[8294]<=26'd11139516; ROM3[8294]<=26'd9750891; ROM4[8294]<=26'd23475089;
ROM1[8295]<=26'd1980510; ROM2[8295]<=26'd11139296; ROM3[8295]<=26'd9753447; ROM4[8295]<=26'd23474811;
ROM1[8296]<=26'd1985524; ROM2[8296]<=26'd11139785; ROM3[8296]<=26'd9753468; ROM4[8296]<=26'd23474878;
ROM1[8297]<=26'd1995334; ROM2[8297]<=26'd11141639; ROM3[8297]<=26'd9751772; ROM4[8297]<=26'd23474104;
ROM1[8298]<=26'd2005181; ROM2[8298]<=26'd11143818; ROM3[8298]<=26'd9746389; ROM4[8298]<=26'd23475524;
ROM1[8299]<=26'd2000925; ROM2[8299]<=26'd11140565; ROM3[8299]<=26'd9740615; ROM4[8299]<=26'd23471645;
ROM1[8300]<=26'd1992023; ROM2[8300]<=26'd11138000; ROM3[8300]<=26'd9739706; ROM4[8300]<=26'd23468433;
ROM1[8301]<=26'd1982484; ROM2[8301]<=26'd11134703; ROM3[8301]<=26'd9739028; ROM4[8301]<=26'd23467168;
ROM1[8302]<=26'd1976747; ROM2[8302]<=26'd11132318; ROM3[8302]<=26'd9739398; ROM4[8302]<=26'd23466491;
ROM1[8303]<=26'd1972897; ROM2[8303]<=26'd11133150; ROM3[8303]<=26'd9742688; ROM4[8303]<=26'd23468247;
ROM1[8304]<=26'd1974375; ROM2[8304]<=26'd11135705; ROM3[8304]<=26'd9744724; ROM4[8304]<=26'd23471741;
ROM1[8305]<=26'd1985233; ROM2[8305]<=26'd11140789; ROM3[8305]<=26'd9745029; ROM4[8305]<=26'd23474898;
ROM1[8306]<=26'd2006306; ROM2[8306]<=26'd11152423; ROM3[8306]<=26'd9749121; ROM4[8306]<=26'd23483988;
ROM1[8307]<=26'd2010675; ROM2[8307]<=26'd11151879; ROM3[8307]<=26'd9745597; ROM4[8307]<=26'd23483711;
ROM1[8308]<=26'd1995383; ROM2[8308]<=26'd11140597; ROM3[8308]<=26'd9736751; ROM4[8308]<=26'd23472645;
ROM1[8309]<=26'd1986451; ROM2[8309]<=26'd11137991; ROM3[8309]<=26'd9738822; ROM4[8309]<=26'd23470790;
ROM1[8310]<=26'd1977216; ROM2[8310]<=26'd11131743; ROM3[8310]<=26'd9739940; ROM4[8310]<=26'd23468254;
ROM1[8311]<=26'd1963114; ROM2[8311]<=26'd11123903; ROM3[8311]<=26'd9735779; ROM4[8311]<=26'd23461114;
ROM1[8312]<=26'd1962755; ROM2[8312]<=26'd11126992; ROM3[8312]<=26'd9737508; ROM4[8312]<=26'd23463083;
ROM1[8313]<=26'd1970080; ROM2[8313]<=26'd11127495; ROM3[8313]<=26'd9736258; ROM4[8313]<=26'd23463538;
ROM1[8314]<=26'd1983370; ROM2[8314]<=26'd11126996; ROM3[8314]<=26'd9730462; ROM4[8314]<=26'd23460458;
ROM1[8315]<=26'd1999195; ROM2[8315]<=26'd11136271; ROM3[8315]<=26'd9732318; ROM4[8315]<=26'd23467359;
ROM1[8316]<=26'd2001670; ROM2[8316]<=26'd11141912; ROM3[8316]<=26'd9740213; ROM4[8316]<=26'd23474037;
ROM1[8317]<=26'd1989723; ROM2[8317]<=26'd11138000; ROM3[8317]<=26'd9740596; ROM4[8317]<=26'd23471806;
ROM1[8318]<=26'd1980101; ROM2[8318]<=26'd11134274; ROM3[8318]<=26'd9738487; ROM4[8318]<=26'd23466899;
ROM1[8319]<=26'd1977703; ROM2[8319]<=26'd11135550; ROM3[8319]<=26'd9742809; ROM4[8319]<=26'd23468600;
ROM1[8320]<=26'd1976728; ROM2[8320]<=26'd11135937; ROM3[8320]<=26'd9742860; ROM4[8320]<=26'd23470179;
ROM1[8321]<=26'd1980820; ROM2[8321]<=26'd11136818; ROM3[8321]<=26'd9739804; ROM4[8321]<=26'd23467889;
ROM1[8322]<=26'd1987137; ROM2[8322]<=26'd11135482; ROM3[8322]<=26'd9732703; ROM4[8322]<=26'd23463902;
ROM1[8323]<=26'd1995059; ROM2[8323]<=26'd11133734; ROM3[8323]<=26'd9726686; ROM4[8323]<=26'd23462365;
ROM1[8324]<=26'd1993462; ROM2[8324]<=26'd11130921; ROM3[8324]<=26'd9725926; ROM4[8324]<=26'd23461285;
ROM1[8325]<=26'd1984893; ROM2[8325]<=26'd11128196; ROM3[8325]<=26'd9727378; ROM4[8325]<=26'd23460699;
ROM1[8326]<=26'd1981627; ROM2[8326]<=26'd11129878; ROM3[8326]<=26'd9732222; ROM4[8326]<=26'd23463338;
ROM1[8327]<=26'd1980516; ROM2[8327]<=26'd11131958; ROM3[8327]<=26'd9737916; ROM4[8327]<=26'd23465274;
ROM1[8328]<=26'd1977771; ROM2[8328]<=26'd11135104; ROM3[8328]<=26'd9743780; ROM4[8328]<=26'd23467824;
ROM1[8329]<=26'd1977583; ROM2[8329]<=26'd11135924; ROM3[8329]<=26'd9743539; ROM4[8329]<=26'd23468257;
ROM1[8330]<=26'd1982741; ROM2[8330]<=26'd11134127; ROM3[8330]<=26'd9737630; ROM4[8330]<=26'd23465841;
ROM1[8331]<=26'd1988457; ROM2[8331]<=26'd11129326; ROM3[8331]<=26'd9726042; ROM4[8331]<=26'd23459276;
ROM1[8332]<=26'd1988579; ROM2[8332]<=26'd11123823; ROM3[8332]<=26'd9717753; ROM4[8332]<=26'd23453656;
ROM1[8333]<=26'd1983666; ROM2[8333]<=26'd11121501; ROM3[8333]<=26'd9718710; ROM4[8333]<=26'd23453342;
ROM1[8334]<=26'd1978372; ROM2[8334]<=26'd11123451; ROM3[8334]<=26'd9725263; ROM4[8334]<=26'd23457124;
ROM1[8335]<=26'd1979624; ROM2[8335]<=26'd11129316; ROM3[8335]<=26'd9733883; ROM4[8335]<=26'd23464075;
ROM1[8336]<=26'd1968704; ROM2[8336]<=26'd11126292; ROM3[8336]<=26'd9735232; ROM4[8336]<=26'd23461816;
ROM1[8337]<=26'd1961109; ROM2[8337]<=26'd11119640; ROM3[8337]<=26'd9729621; ROM4[8337]<=26'd23455388;
ROM1[8338]<=26'd1965701; ROM2[8338]<=26'd11117972; ROM3[8338]<=26'd9723996; ROM4[8338]<=26'd23453037;
ROM1[8339]<=26'd1977276; ROM2[8339]<=26'd11117816; ROM3[8339]<=26'd9720992; ROM4[8339]<=26'd23454141;
ROM1[8340]<=26'd1989786; ROM2[8340]<=26'd11122314; ROM3[8340]<=26'd9721564; ROM4[8340]<=26'd23458267;
ROM1[8341]<=26'd1996597; ROM2[8341]<=26'd11134592; ROM3[8341]<=26'd9734982; ROM4[8341]<=26'd23469729;
ROM1[8342]<=26'd1987746; ROM2[8342]<=26'd11133439; ROM3[8342]<=26'd9739747; ROM4[8342]<=26'd23471011;
ROM1[8343]<=26'd1973738; ROM2[8343]<=26'd11124532; ROM3[8343]<=26'd9733895; ROM4[8343]<=26'd23462697;
ROM1[8344]<=26'd1965556; ROM2[8344]<=26'd11121100; ROM3[8344]<=26'd9734190; ROM4[8344]<=26'd23459761;
ROM1[8345]<=26'd1956540; ROM2[8345]<=26'd11114384; ROM3[8345]<=26'd9732123; ROM4[8345]<=26'd23455294;
ROM1[8346]<=26'd1957623; ROM2[8346]<=26'd11114817; ROM3[8346]<=26'd9729416; ROM4[8346]<=26'd23453339;
ROM1[8347]<=26'd1972919; ROM2[8347]<=26'd11121585; ROM3[8347]<=26'd9729707; ROM4[8347]<=26'd23457545;
ROM1[8348]<=26'd1986692; ROM2[8348]<=26'd11124027; ROM3[8348]<=26'd9725655; ROM4[8348]<=26'd23458709;
ROM1[8349]<=26'd1989402; ROM2[8349]<=26'd11127825; ROM3[8349]<=26'd9726363; ROM4[8349]<=26'd23461200;
ROM1[8350]<=26'd1993403; ROM2[8350]<=26'd11136489; ROM3[8350]<=26'd9739278; ROM4[8350]<=26'd23471292;
ROM1[8351]<=26'd1982878; ROM2[8351]<=26'd11132919; ROM3[8351]<=26'd9739819; ROM4[8351]<=26'd23469202;
ROM1[8352]<=26'd1967103; ROM2[8352]<=26'd11122088; ROM3[8352]<=26'd9732370; ROM4[8352]<=26'd23460131;
ROM1[8353]<=26'd1960562; ROM2[8353]<=26'd11119034; ROM3[8353]<=26'd9731480; ROM4[8353]<=26'd23457043;
ROM1[8354]<=26'd1955601; ROM2[8354]<=26'd11112240; ROM3[8354]<=26'd9722834; ROM4[8354]<=26'd23450184;
ROM1[8355]<=26'd1965797; ROM2[8355]<=26'd11114149; ROM3[8355]<=26'd9721148; ROM4[8355]<=26'd23450975;
ROM1[8356]<=26'd1986264; ROM2[8356]<=26'd11123026; ROM3[8356]<=26'd9725044; ROM4[8356]<=26'd23458811;
ROM1[8357]<=26'd1987967; ROM2[8357]<=26'd11120103; ROM3[8357]<=26'd9722648; ROM4[8357]<=26'd23457765;
ROM1[8358]<=26'd1982503; ROM2[8358]<=26'd11118825; ROM3[8358]<=26'd9725166; ROM4[8358]<=26'd23455675;
ROM1[8359]<=26'd1982191; ROM2[8359]<=26'd11124107; ROM3[8359]<=26'd9735206; ROM4[8359]<=26'd23462338;
ROM1[8360]<=26'd1977962; ROM2[8360]<=26'd11124389; ROM3[8360]<=26'd9737279; ROM4[8360]<=26'd23462899;
ROM1[8361]<=26'd1966189; ROM2[8361]<=26'd11118846; ROM3[8361]<=26'd9732819; ROM4[8361]<=26'd23456120;
ROM1[8362]<=26'd1968818; ROM2[8362]<=26'd11123297; ROM3[8362]<=26'd9738681; ROM4[8362]<=26'd23462309;
ROM1[8363]<=26'd1975930; ROM2[8363]<=26'd11125717; ROM3[8363]<=26'd9737415; ROM4[8363]<=26'd23463105;
ROM1[8364]<=26'd1984949; ROM2[8364]<=26'd11124805; ROM3[8364]<=26'd9731075; ROM4[8364]<=26'd23459371;
ROM1[8365]<=26'd1995148; ROM2[8365]<=26'd11126216; ROM3[8365]<=26'd9728433; ROM4[8365]<=26'd23461554;
ROM1[8366]<=26'd1992124; ROM2[8366]<=26'd11125435; ROM3[8366]<=26'd9729676; ROM4[8366]<=26'd23460753;
ROM1[8367]<=26'd1985225; ROM2[8367]<=26'd11126184; ROM3[8367]<=26'd9733443; ROM4[8367]<=26'd23460832;
ROM1[8368]<=26'd1977901; ROM2[8368]<=26'd11125246; ROM3[8368]<=26'd9734522; ROM4[8368]<=26'd23460872;
ROM1[8369]<=26'd1972457; ROM2[8369]<=26'd11125612; ROM3[8369]<=26'd9737357; ROM4[8369]<=26'd23459800;
ROM1[8370]<=26'd1960284; ROM2[8370]<=26'd11118208; ROM3[8370]<=26'd9728891; ROM4[8370]<=26'd23451528;
ROM1[8371]<=26'd1957652; ROM2[8371]<=26'd11113491; ROM3[8371]<=26'd9722236; ROM4[8371]<=26'd23446598;
ROM1[8372]<=26'd1971809; ROM2[8372]<=26'd11117809; ROM3[8372]<=26'd9721224; ROM4[8372]<=26'd23447386;
ROM1[8373]<=26'd1982666; ROM2[8373]<=26'd11120302; ROM3[8373]<=26'd9717206; ROM4[8373]<=26'd23447641;
ROM1[8374]<=26'd1979743; ROM2[8374]<=26'd11118207; ROM3[8374]<=26'd9716923; ROM4[8374]<=26'd23447237;
ROM1[8375]<=26'd1974591; ROM2[8375]<=26'd11118119; ROM3[8375]<=26'd9721659; ROM4[8375]<=26'd23449625;
ROM1[8376]<=26'd1975611; ROM2[8376]<=26'd11125675; ROM3[8376]<=26'd9732214; ROM4[8376]<=26'd23458551;
ROM1[8377]<=26'd1970094; ROM2[8377]<=26'd11125624; ROM3[8377]<=26'd9733309; ROM4[8377]<=26'd23458777;
ROM1[8378]<=26'd1962901; ROM2[8378]<=26'd11123059; ROM3[8378]<=26'd9733457; ROM4[8378]<=26'd23457146;
ROM1[8379]<=26'd1960026; ROM2[8379]<=26'd11120132; ROM3[8379]<=26'd9730381; ROM4[8379]<=26'd23454218;
ROM1[8380]<=26'd1960249; ROM2[8380]<=26'd11112637; ROM3[8380]<=26'd9720153; ROM4[8380]<=26'd23446395;
ROM1[8381]<=26'd1971346; ROM2[8381]<=26'd11113177; ROM3[8381]<=26'd9714215; ROM4[8381]<=26'd23445855;
ROM1[8382]<=26'd1978135; ROM2[8382]<=26'd11118001; ROM3[8382]<=26'd9715605; ROM4[8382]<=26'd23449786;
ROM1[8383]<=26'd1973283; ROM2[8383]<=26'd11117434; ROM3[8383]<=26'd9717025; ROM4[8383]<=26'd23449321;
ROM1[8384]<=26'd1967667; ROM2[8384]<=26'd11117270; ROM3[8384]<=26'd9720793; ROM4[8384]<=26'd23451502;
ROM1[8385]<=26'd1965384; ROM2[8385]<=26'd11117953; ROM3[8385]<=26'd9726250; ROM4[8385]<=26'd23453738;
ROM1[8386]<=26'd1959442; ROM2[8386]<=26'd11117010; ROM3[8386]<=26'd9727267; ROM4[8386]<=26'd23451950;
ROM1[8387]<=26'd1957667; ROM2[8387]<=26'd11117610; ROM3[8387]<=26'd9726567; ROM4[8387]<=26'd23451427;
ROM1[8388]<=26'd1962965; ROM2[8388]<=26'd11118951; ROM3[8388]<=26'd9726197; ROM4[8388]<=26'd23451168;
ROM1[8389]<=26'd1978133; ROM2[8389]<=26'd11123877; ROM3[8389]<=26'd9722941; ROM4[8389]<=26'd23453325;
ROM1[8390]<=26'd1987319; ROM2[8390]<=26'd11125486; ROM3[8390]<=26'd9718807; ROM4[8390]<=26'd23452432;
ROM1[8391]<=26'd1984902; ROM2[8391]<=26'd11125821; ROM3[8391]<=26'd9721509; ROM4[8391]<=26'd23452894;
ROM1[8392]<=26'd1975765; ROM2[8392]<=26'd11124196; ROM3[8392]<=26'd9721935; ROM4[8392]<=26'd23451008;
ROM1[8393]<=26'd1968014; ROM2[8393]<=26'd11122047; ROM3[8393]<=26'd9725066; ROM4[8393]<=26'd23450864;
ROM1[8394]<=26'd1961039; ROM2[8394]<=26'd11121235; ROM3[8394]<=26'd9727509; ROM4[8394]<=26'd23450305;
ROM1[8395]<=26'd1957664; ROM2[8395]<=26'd11122581; ROM3[8395]<=26'd9730313; ROM4[8395]<=26'd23450206;
ROM1[8396]<=26'd1968270; ROM2[8396]<=26'd11132098; ROM3[8396]<=26'd9739330; ROM4[8396]<=26'd23459570;
ROM1[8397]<=26'd1982693; ROM2[8397]<=26'd11136854; ROM3[8397]<=26'd9740671; ROM4[8397]<=26'd23464438;
ROM1[8398]<=26'd1988397; ROM2[8398]<=26'd11130757; ROM3[8398]<=26'd9730607; ROM4[8398]<=26'd23459874;
ROM1[8399]<=26'd1981049; ROM2[8399]<=26'd11123990; ROM3[8399]<=26'd9723952; ROM4[8399]<=26'd23455272;
ROM1[8400]<=26'd1974079; ROM2[8400]<=26'd11122352; ROM3[8400]<=26'd9726900; ROM4[8400]<=26'd23454314;
ROM1[8401]<=26'd1970827; ROM2[8401]<=26'd11123992; ROM3[8401]<=26'd9732688; ROM4[8401]<=26'd23457371;
ROM1[8402]<=26'd1969676; ROM2[8402]<=26'd11128325; ROM3[8402]<=26'd9738800; ROM4[8402]<=26'd23463009;
ROM1[8403]<=26'd1971586; ROM2[8403]<=26'd11135448; ROM3[8403]<=26'd9748436; ROM4[8403]<=26'd23470285;
ROM1[8404]<=26'd1978810; ROM2[8404]<=26'd11140733; ROM3[8404]<=26'd9752768; ROM4[8404]<=26'd23476627;
ROM1[8405]<=26'd1978934; ROM2[8405]<=26'd11132527; ROM3[8405]<=26'd9740413; ROM4[8405]<=26'd23467572;
ROM1[8406]<=26'd1986724; ROM2[8406]<=26'd11127217; ROM3[8406]<=26'd9729237; ROM4[8406]<=26'd23460199;
ROM1[8407]<=26'd1990882; ROM2[8407]<=26'd11126401; ROM3[8407]<=26'd9726834; ROM4[8407]<=26'd23459442;
ROM1[8408]<=26'd1981554; ROM2[8408]<=26'd11123429; ROM3[8408]<=26'd9725794; ROM4[8408]<=26'd23456907;
ROM1[8409]<=26'd1976099; ROM2[8409]<=26'd11125800; ROM3[8409]<=26'd9733237; ROM4[8409]<=26'd23461613;
ROM1[8410]<=26'd1975301; ROM2[8410]<=26'd11129015; ROM3[8410]<=26'd9741576; ROM4[8410]<=26'd23467522;
ROM1[8411]<=26'd1967136; ROM2[8411]<=26'd11124904; ROM3[8411]<=26'd9742424; ROM4[8411]<=26'd23465289;
ROM1[8412]<=26'd1962046; ROM2[8412]<=26'd11121026; ROM3[8412]<=26'd9737378; ROM4[8412]<=26'd23460073;
ROM1[8413]<=26'd1968494; ROM2[8413]<=26'd11121339; ROM3[8413]<=26'd9733210; ROM4[8413]<=26'd23457414;
ROM1[8414]<=26'd1978258; ROM2[8414]<=26'd11121608; ROM3[8414]<=26'd9727819; ROM4[8414]<=26'd23456073;
ROM1[8415]<=26'd1981977; ROM2[8415]<=26'd11120199; ROM3[8415]<=26'd9720153; ROM4[8415]<=26'd23454731;
ROM1[8416]<=26'd1973302; ROM2[8416]<=26'd11114527; ROM3[8416]<=26'd9717881; ROM4[8416]<=26'd23450510;
ROM1[8417]<=26'd1962949; ROM2[8417]<=26'd11112162; ROM3[8417]<=26'd9719792; ROM4[8417]<=26'd23448791;
ROM1[8418]<=26'd1960390; ROM2[8418]<=26'd11114159; ROM3[8418]<=26'd9723014; ROM4[8418]<=26'd23451128;
ROM1[8419]<=26'd1954222; ROM2[8419]<=26'd11113457; ROM3[8419]<=26'd9724238; ROM4[8419]<=26'd23450046;
ROM1[8420]<=26'd1949453; ROM2[8420]<=26'd11111703; ROM3[8420]<=26'd9722660; ROM4[8420]<=26'd23447568;
ROM1[8421]<=26'd1953280; ROM2[8421]<=26'd11113293; ROM3[8421]<=26'd9720511; ROM4[8421]<=26'd23446616;
ROM1[8422]<=26'd1962668; ROM2[8422]<=26'd11115633; ROM3[8422]<=26'd9717521; ROM4[8422]<=26'd23446277;
ROM1[8423]<=26'd1974068; ROM2[8423]<=26'd11116066; ROM3[8423]<=26'd9712628; ROM4[8423]<=26'd23445088;
ROM1[8424]<=26'd1972330; ROM2[8424]<=26'd11115714; ROM3[8424]<=26'd9711918; ROM4[8424]<=26'd23443782;
ROM1[8425]<=26'd1963221; ROM2[8425]<=26'd11113755; ROM3[8425]<=26'd9712598; ROM4[8425]<=26'd23442440;
ROM1[8426]<=26'd1958031; ROM2[8426]<=26'd11111453; ROM3[8426]<=26'd9713857; ROM4[8426]<=26'd23442445;
ROM1[8427]<=26'd1953199; ROM2[8427]<=26'd11110369; ROM3[8427]<=26'd9714253; ROM4[8427]<=26'd23441274;
ROM1[8428]<=26'd1946291; ROM2[8428]<=26'd11108141; ROM3[8428]<=26'd9714177; ROM4[8428]<=26'd23439439;
ROM1[8429]<=26'd1947586; ROM2[8429]<=26'd11107661; ROM3[8429]<=26'd9714302; ROM4[8429]<=26'd23439145;
ROM1[8430]<=26'd1955003; ROM2[8430]<=26'd11110850; ROM3[8430]<=26'd9712343; ROM4[8430]<=26'd23440213;
ROM1[8431]<=26'd1965829; ROM2[8431]<=26'd11111537; ROM3[8431]<=26'd9706379; ROM4[8431]<=26'd23439662;
ROM1[8432]<=26'd1970421; ROM2[8432]<=26'd11112193; ROM3[8432]<=26'd9705079; ROM4[8432]<=26'd23440696;
ROM1[8433]<=26'd1968483; ROM2[8433]<=26'd11114407; ROM3[8433]<=26'd9711299; ROM4[8433]<=26'd23445768;
ROM1[8434]<=26'd1961884; ROM2[8434]<=26'd11111444; ROM3[8434]<=26'd9714081; ROM4[8434]<=26'd23444003;
ROM1[8435]<=26'd1953761; ROM2[8435]<=26'd11106527; ROM3[8435]<=26'd9715687; ROM4[8435]<=26'd23441079;
ROM1[8436]<=26'd1945031; ROM2[8436]<=26'd11103980; ROM3[8436]<=26'd9716362; ROM4[8436]<=26'd23440168;
ROM1[8437]<=26'd1942789; ROM2[8437]<=26'd11104440; ROM3[8437]<=26'd9715435; ROM4[8437]<=26'd23439961;
ROM1[8438]<=26'd1951443; ROM2[8438]<=26'd11107126; ROM3[8438]<=26'd9716615; ROM4[8438]<=26'd23443278;
ROM1[8439]<=26'd1973180; ROM2[8439]<=26'd11116444; ROM3[8439]<=26'd9721584; ROM4[8439]<=26'd23452882;
ROM1[8440]<=26'd1988667; ROM2[8440]<=26'd11121618; ROM3[8440]<=26'd9727906; ROM4[8440]<=26'd23462593;
ROM1[8441]<=26'd1976462; ROM2[8441]<=26'd11110862; ROM3[8441]<=26'd9721909; ROM4[8441]<=26'd23455734;
ROM1[8442]<=26'd1969127; ROM2[8442]<=26'd11111552; ROM3[8442]<=26'd9727406; ROM4[8442]<=26'd23456544;
ROM1[8443]<=26'd1970255; ROM2[8443]<=26'd11119593; ROM3[8443]<=26'd9738047; ROM4[8443]<=26'd23464307;
ROM1[8444]<=26'd1962131; ROM2[8444]<=26'd11115704; ROM3[8444]<=26'd9732547; ROM4[8444]<=26'd23458864;
ROM1[8445]<=26'd1964869; ROM2[8445]<=26'd11122301; ROM3[8445]<=26'd9734944; ROM4[8445]<=26'd23461225;
ROM1[8446]<=26'd1967554; ROM2[8446]<=26'd11121673; ROM3[8446]<=26'd9730230; ROM4[8446]<=26'd23457261;
ROM1[8447]<=26'd1970537; ROM2[8447]<=26'd11113311; ROM3[8447]<=26'd9719966; ROM4[8447]<=26'd23448762;
ROM1[8448]<=26'd1982541; ROM2[8448]<=26'd11116882; ROM3[8448]<=26'd9717792; ROM4[8448]<=26'd23450775;
ROM1[8449]<=26'd1980977; ROM2[8449]<=26'd11116872; ROM3[8449]<=26'd9718521; ROM4[8449]<=26'd23450983;
ROM1[8450]<=26'd1973588; ROM2[8450]<=26'd11115233; ROM3[8450]<=26'd9721260; ROM4[8450]<=26'd23450362;
ROM1[8451]<=26'd1976731; ROM2[8451]<=26'd11123135; ROM3[8451]<=26'd9729316; ROM4[8451]<=26'd23457269;
ROM1[8452]<=26'd1975362; ROM2[8452]<=26'd11126187; ROM3[8452]<=26'd9734655; ROM4[8452]<=26'd23460557;
ROM1[8453]<=26'd1967347; ROM2[8453]<=26'd11121726; ROM3[8453]<=26'd9735730; ROM4[8453]<=26'd23456666;
ROM1[8454]<=26'd1967810; ROM2[8454]<=26'd11120276; ROM3[8454]<=26'd9734605; ROM4[8454]<=26'd23456011;
ROM1[8455]<=26'd1974160; ROM2[8455]<=26'd11122544; ROM3[8455]<=26'd9728301; ROM4[8455]<=26'd23455533;
ROM1[8456]<=26'd1984017; ROM2[8456]<=26'd11121416; ROM3[8456]<=26'd9721352; ROM4[8456]<=26'd23451270;
ROM1[8457]<=26'd1988515; ROM2[8457]<=26'd11119786; ROM3[8457]<=26'd9720224; ROM4[8457]<=26'd23450896;
ROM1[8458]<=26'd1983333; ROM2[8458]<=26'd11120158; ROM3[8458]<=26'd9722658; ROM4[8458]<=26'd23453419;
ROM1[8459]<=26'd1971627; ROM2[8459]<=26'd11114023; ROM3[8459]<=26'd9724906; ROM4[8459]<=26'd23450416;
ROM1[8460]<=26'd1964894; ROM2[8460]<=26'd11114144; ROM3[8460]<=26'd9727640; ROM4[8460]<=26'd23451052;
ROM1[8461]<=26'd1962482; ROM2[8461]<=26'd11118652; ROM3[8461]<=26'd9732700; ROM4[8461]<=26'd23456140;
ROM1[8462]<=26'd1960277; ROM2[8462]<=26'd11117996; ROM3[8462]<=26'd9734332; ROM4[8462]<=26'd23457446;
ROM1[8463]<=26'd1961690; ROM2[8463]<=26'd11115184; ROM3[8463]<=26'd9728663; ROM4[8463]<=26'd23455048;
ROM1[8464]<=26'd1974024; ROM2[8464]<=26'd11117208; ROM3[8464]<=26'd9723926; ROM4[8464]<=26'd23454763;
ROM1[8465]<=26'd1982941; ROM2[8465]<=26'd11122223; ROM3[8465]<=26'd9721197; ROM4[8465]<=26'd23457835;
ROM1[8466]<=26'd1978103; ROM2[8466]<=26'd11122077; ROM3[8466]<=26'd9720119; ROM4[8466]<=26'd23458970;
ROM1[8467]<=26'd1968698; ROM2[8467]<=26'd11120461; ROM3[8467]<=26'd9720238; ROM4[8467]<=26'd23457142;
ROM1[8468]<=26'd1962472; ROM2[8468]<=26'd11118984; ROM3[8468]<=26'd9720740; ROM4[8468]<=26'd23456155;
ROM1[8469]<=26'd1954016; ROM2[8469]<=26'd11114864; ROM3[8469]<=26'd9720809; ROM4[8469]<=26'd23453123;
ROM1[8470]<=26'd1948804; ROM2[8470]<=26'd11115064; ROM3[8470]<=26'd9721252; ROM4[8470]<=26'd23451974;
ROM1[8471]<=26'd1952939; ROM2[8471]<=26'd11118005; ROM3[8471]<=26'd9719842; ROM4[8471]<=26'd23451659;
ROM1[8472]<=26'd1966512; ROM2[8472]<=26'd11121815; ROM3[8472]<=26'd9717250; ROM4[8472]<=26'd23453926;
ROM1[8473]<=26'd1979798; ROM2[8473]<=26'd11125355; ROM3[8473]<=26'd9714736; ROM4[8473]<=26'd23456368;
ROM1[8474]<=26'd1975641; ROM2[8474]<=26'd11121986; ROM3[8474]<=26'd9710681; ROM4[8474]<=26'd23451677;
ROM1[8475]<=26'd1966676; ROM2[8475]<=26'd11119044; ROM3[8475]<=26'd9709765; ROM4[8475]<=26'd23447403;
ROM1[8476]<=26'd1956989; ROM2[8476]<=26'd11116368; ROM3[8476]<=26'd9710224; ROM4[8476]<=26'd23442929;
ROM1[8477]<=26'd1950015; ROM2[8477]<=26'd11113036; ROM3[8477]<=26'd9710522; ROM4[8477]<=26'd23439509;
ROM1[8478]<=26'd1946152; ROM2[8478]<=26'd11113275; ROM3[8478]<=26'd9712621; ROM4[8478]<=26'd23439847;
ROM1[8479]<=26'd1949451; ROM2[8479]<=26'd11115259; ROM3[8479]<=26'd9716716; ROM4[8479]<=26'd23442145;
ROM1[8480]<=26'd1959303; ROM2[8480]<=26'd11116186; ROM3[8480]<=26'd9716207; ROM4[8480]<=26'd23442851;
ROM1[8481]<=26'd1972627; ROM2[8481]<=26'd11118568; ROM3[8481]<=26'd9710550; ROM4[8481]<=26'd23443775;
ROM1[8482]<=26'd1973616; ROM2[8482]<=26'd11116985; ROM3[8482]<=26'd9708596; ROM4[8482]<=26'd23441320;
ROM1[8483]<=26'd1960886; ROM2[8483]<=26'd11108352; ROM3[8483]<=26'd9705973; ROM4[8483]<=26'd23435210;
ROM1[8484]<=26'd1958694; ROM2[8484]<=26'd11112311; ROM3[8484]<=26'd9713947; ROM4[8484]<=26'd23441091;
ROM1[8485]<=26'd1955223; ROM2[8485]<=26'd11115315; ROM3[8485]<=26'd9719346; ROM4[8485]<=26'd23443313;
ROM1[8486]<=26'd1943822; ROM2[8486]<=26'd11108168; ROM3[8486]<=26'd9714726; ROM4[8486]<=26'd23436001;
ROM1[8487]<=26'd1946487; ROM2[8487]<=26'd11111790; ROM3[8487]<=26'd9716567; ROM4[8487]<=26'd23438133;
ROM1[8488]<=26'd1952113; ROM2[8488]<=26'd11111587; ROM3[8488]<=26'd9714215; ROM4[8488]<=26'd23437941;
ROM1[8489]<=26'd1964499; ROM2[8489]<=26'd11112618; ROM3[8489]<=26'd9709637; ROM4[8489]<=26'd23437864;
ROM1[8490]<=26'd1979458; ROM2[8490]<=26'd11121689; ROM3[8490]<=26'd9712814; ROM4[8490]<=26'd23446003;
ROM1[8491]<=26'd1970517; ROM2[8491]<=26'd11117380; ROM3[8491]<=26'd9709346; ROM4[8491]<=26'd23443911;
ROM1[8492]<=26'd1957552; ROM2[8492]<=26'd11112740; ROM3[8492]<=26'd9707141; ROM4[8492]<=26'd23439501;
ROM1[8493]<=26'd1948042; ROM2[8493]<=26'd11108976; ROM3[8493]<=26'd9706901; ROM4[8493]<=26'd23436651;
ROM1[8494]<=26'd1944443; ROM2[8494]<=26'd11108323; ROM3[8494]<=26'd9710487; ROM4[8494]<=26'd23438784;
ROM1[8495]<=26'd1948080; ROM2[8495]<=26'd11112414; ROM3[8495]<=26'd9716070; ROM4[8495]<=26'd23444008;
ROM1[8496]<=26'd1951969; ROM2[8496]<=26'd11112883; ROM3[8496]<=26'd9715181; ROM4[8496]<=26'd23443677;
ROM1[8497]<=26'd1964096; ROM2[8497]<=26'd11115325; ROM3[8497]<=26'd9713399; ROM4[8497]<=26'd23444636;
ROM1[8498]<=26'd1977804; ROM2[8498]<=26'd11118010; ROM3[8498]<=26'd9709647; ROM4[8498]<=26'd23444755;
ROM1[8499]<=26'd1980264; ROM2[8499]<=26'd11121576; ROM3[8499]<=26'd9711306; ROM4[8499]<=26'd23449021;
ROM1[8500]<=26'd1972953; ROM2[8500]<=26'd11122729; ROM3[8500]<=26'd9714128; ROM4[8500]<=26'd23450403;
ROM1[8501]<=26'd1970746; ROM2[8501]<=26'd11125939; ROM3[8501]<=26'd9720818; ROM4[8501]<=26'd23452736;
ROM1[8502]<=26'd1969957; ROM2[8502]<=26'd11127906; ROM3[8502]<=26'd9727856; ROM4[8502]<=26'd23457874;
ROM1[8503]<=26'd1955124; ROM2[8503]<=26'd11116911; ROM3[8503]<=26'd9721749; ROM4[8503]<=26'd23449036;
ROM1[8504]<=26'd1952664; ROM2[8504]<=26'd11112372; ROM3[8504]<=26'd9716348; ROM4[8504]<=26'd23443563;
ROM1[8505]<=26'd1963969; ROM2[8505]<=26'd11116654; ROM3[8505]<=26'd9714267; ROM4[8505]<=26'd23445120;
ROM1[8506]<=26'd1975320; ROM2[8506]<=26'd11119224; ROM3[8506]<=26'd9709465; ROM4[8506]<=26'd23443317;
ROM1[8507]<=26'd1980223; ROM2[8507]<=26'd11123674; ROM3[8507]<=26'd9710759; ROM4[8507]<=26'd23445165;
ROM1[8508]<=26'd1973885; ROM2[8508]<=26'd11121834; ROM3[8508]<=26'd9712447; ROM4[8508]<=26'd23445551;
ROM1[8509]<=26'd1967274; ROM2[8509]<=26'd11120071; ROM3[8509]<=26'd9717416; ROM4[8509]<=26'd23447881;
ROM1[8510]<=26'd1960337; ROM2[8510]<=26'd11118336; ROM3[8510]<=26'd9720235; ROM4[8510]<=26'd23447649;
ROM1[8511]<=26'd1959393; ROM2[8511]<=26'd11121826; ROM3[8511]<=26'd9728523; ROM4[8511]<=26'd23452192;
ROM1[8512]<=26'd1962279; ROM2[8512]<=26'd11127000; ROM3[8512]<=26'd9732771; ROM4[8512]<=26'd23456619;
ROM1[8513]<=26'd1962351; ROM2[8513]<=26'd11122181; ROM3[8513]<=26'd9723680; ROM4[8513]<=26'd23450880;
ROM1[8514]<=26'd1970866; ROM2[8514]<=26'd11118656; ROM3[8514]<=26'd9714269; ROM4[8514]<=26'd23446661;
ROM1[8515]<=26'd1975562; ROM2[8515]<=26'd11115773; ROM3[8515]<=26'd9707230; ROM4[8515]<=26'd23442054;
ROM1[8516]<=26'd1973837; ROM2[8516]<=26'd11114911; ROM3[8516]<=26'd9708135; ROM4[8516]<=26'd23441328;
ROM1[8517]<=26'd1968009; ROM2[8517]<=26'd11114057; ROM3[8517]<=26'd9712044; ROM4[8517]<=26'd23441007;
ROM1[8518]<=26'd1958788; ROM2[8518]<=26'd11113284; ROM3[8518]<=26'd9712022; ROM4[8518]<=26'd23439214;
ROM1[8519]<=26'd1954516; ROM2[8519]<=26'd11114708; ROM3[8519]<=26'd9715116; ROM4[8519]<=26'd23440377;
ROM1[8520]<=26'd1950044; ROM2[8520]<=26'd11112982; ROM3[8520]<=26'd9715619; ROM4[8520]<=26'd23439741;
ROM1[8521]<=26'd1949408; ROM2[8521]<=26'd11110690; ROM3[8521]<=26'd9709619; ROM4[8521]<=26'd23435192;
ROM1[8522]<=26'd1958256; ROM2[8522]<=26'd11108691; ROM3[8522]<=26'd9701827; ROM4[8522]<=26'd23431238;
ROM1[8523]<=26'd1973421; ROM2[8523]<=26'd11114876; ROM3[8523]<=26'd9701194; ROM4[8523]<=26'd23436177;
ROM1[8524]<=26'd1968135; ROM2[8524]<=26'd11112198; ROM3[8524]<=26'd9700251; ROM4[8524]<=26'd23433907;
ROM1[8525]<=26'd1952548; ROM2[8525]<=26'd11101903; ROM3[8525]<=26'd9696564; ROM4[8525]<=26'd23428160;
ROM1[8526]<=26'd1947278; ROM2[8526]<=26'd11102930; ROM3[8526]<=26'd9701916; ROM4[8526]<=26'd23430237;
ROM1[8527]<=26'd1939665; ROM2[8527]<=26'd11100021; ROM3[8527]<=26'd9701682; ROM4[8527]<=26'd23428655;
ROM1[8528]<=26'd1932333; ROM2[8528]<=26'd11096517; ROM3[8528]<=26'd9700509; ROM4[8528]<=26'd23426579;
ROM1[8529]<=26'd1935863; ROM2[8529]<=26'd11099782; ROM3[8529]<=26'd9703114; ROM4[8529]<=26'd23428502;
ROM1[8530]<=26'd1949601; ROM2[8530]<=26'd11105482; ROM3[8530]<=26'd9705569; ROM4[8530]<=26'd23433449;
ROM1[8531]<=26'd1964988; ROM2[8531]<=26'd11109216; ROM3[8531]<=26'd9704092; ROM4[8531]<=26'd23437976;
ROM1[8532]<=26'd1971662; ROM2[8532]<=26'd11111798; ROM3[8532]<=26'd9707479; ROM4[8532]<=26'd23442942;
ROM1[8533]<=26'd1971481; ROM2[8533]<=26'd11116751; ROM3[8533]<=26'd9716959; ROM4[8533]<=26'd23449325;
ROM1[8534]<=26'd1963111; ROM2[8534]<=26'd11116601; ROM3[8534]<=26'd9720589; ROM4[8534]<=26'd23449857;
ROM1[8535]<=26'd1950847; ROM2[8535]<=26'd11109926; ROM3[8535]<=26'd9716108; ROM4[8535]<=26'd23440771;
ROM1[8536]<=26'd1940677; ROM2[8536]<=26'd11104430; ROM3[8536]<=26'd9712717; ROM4[8536]<=26'd23434759;
ROM1[8537]<=26'd1936301; ROM2[8537]<=26'd11100067; ROM3[8537]<=26'd9708394; ROM4[8537]<=26'd23430781;
ROM1[8538]<=26'd1939686; ROM2[8538]<=26'd11097825; ROM3[8538]<=26'd9702406; ROM4[8538]<=26'd23427468;
ROM1[8539]<=26'd1955172; ROM2[8539]<=26'd11102319; ROM3[8539]<=26'd9699824; ROM4[8539]<=26'd23429894;
ROM1[8540]<=26'd1964828; ROM2[8540]<=26'd11106565; ROM3[8540]<=26'd9698083; ROM4[8540]<=26'd23432870;
ROM1[8541]<=26'd1960497; ROM2[8541]<=26'd11106683; ROM3[8541]<=26'd9698138; ROM4[8541]<=26'd23433877;
ROM1[8542]<=26'd1955588; ROM2[8542]<=26'd11105295; ROM3[8542]<=26'd9702178; ROM4[8542]<=26'd23435040;
ROM1[8543]<=26'd1951311; ROM2[8543]<=26'd11105590; ROM3[8543]<=26'd9707973; ROM4[8543]<=26'd23437701;
ROM1[8544]<=26'd1949393; ROM2[8544]<=26'd11111205; ROM3[8544]<=26'd9717140; ROM4[8544]<=26'd23443721;
ROM1[8545]<=26'd1948959; ROM2[8545]<=26'd11112640; ROM3[8545]<=26'd9721382; ROM4[8545]<=26'd23445726;
ROM1[8546]<=26'd1950587; ROM2[8546]<=26'd11109939; ROM3[8546]<=26'd9715741; ROM4[8546]<=26'd23442734;
ROM1[8547]<=26'd1963116; ROM2[8547]<=26'd11112181; ROM3[8547]<=26'd9711864; ROM4[8547]<=26'd23445024;
ROM1[8548]<=26'd1979876; ROM2[8548]<=26'd11116994; ROM3[8548]<=26'd9713258; ROM4[8548]<=26'd23451102;
ROM1[8549]<=26'd1978074; ROM2[8549]<=26'd11117212; ROM3[8549]<=26'd9713077; ROM4[8549]<=26'd23452421;
ROM1[8550]<=26'd1963047; ROM2[8550]<=26'd11110556; ROM3[8550]<=26'd9707640; ROM4[8550]<=26'd23445528;
ROM1[8551]<=26'd1953004; ROM2[8551]<=26'd11105293; ROM3[8551]<=26'd9706459; ROM4[8551]<=26'd23439104;
ROM1[8552]<=26'd1946399; ROM2[8552]<=26'd11101952; ROM3[8552]<=26'd9704851; ROM4[8552]<=26'd23436605;
ROM1[8553]<=26'd1939354; ROM2[8553]<=26'd11100254; ROM3[8553]<=26'd9705385; ROM4[8553]<=26'd23434871;
ROM1[8554]<=26'd1947110; ROM2[8554]<=26'd11106708; ROM3[8554]<=26'd9711556; ROM4[8554]<=26'd23439474;
ROM1[8555]<=26'd1956803; ROM2[8555]<=26'd11108968; ROM3[8555]<=26'd9706826; ROM4[8555]<=26'd23438976;
ROM1[8556]<=26'd1967996; ROM2[8556]<=26'd11109120; ROM3[8556]<=26'd9698922; ROM4[8556]<=26'd23436338;
ROM1[8557]<=26'd1975587; ROM2[8557]<=26'd11113148; ROM3[8557]<=26'd9699515; ROM4[8557]<=26'd23439877;
ROM1[8558]<=26'd1973735; ROM2[8558]<=26'd11117644; ROM3[8558]<=26'd9706679; ROM4[8558]<=26'd23445121;
ROM1[8559]<=26'd1971915; ROM2[8559]<=26'd11126229; ROM3[8559]<=26'd9718567; ROM4[8559]<=26'd23453886;
ROM1[8560]<=26'd1966245; ROM2[8560]<=26'd11127749; ROM3[8560]<=26'd9722108; ROM4[8560]<=26'd23454981;
ROM1[8561]<=26'd1950892; ROM2[8561]<=26'd11117611; ROM3[8561]<=26'd9716620; ROM4[8561]<=26'd23444216;
ROM1[8562]<=26'd1944030; ROM2[8562]<=26'd11112383; ROM3[8562]<=26'd9710228; ROM4[8562]<=26'd23439144;
ROM1[8563]<=26'd1951093; ROM2[8563]<=26'd11112239; ROM3[8563]<=26'd9706235; ROM4[8563]<=26'd23439966;
ROM1[8564]<=26'd1964305; ROM2[8564]<=26'd11113159; ROM3[8564]<=26'd9700801; ROM4[8564]<=26'd23438690;
ROM1[8565]<=26'd1978222; ROM2[8565]<=26'd11122430; ROM3[8565]<=26'd9703344; ROM4[8565]<=26'd23445438;
ROM1[8566]<=26'd1976693; ROM2[8566]<=26'd11125581; ROM3[8566]<=26'd9708184; ROM4[8566]<=26'd23449021;
ROM1[8567]<=26'd1959221; ROM2[8567]<=26'd11113715; ROM3[8567]<=26'd9701799; ROM4[8567]<=26'd23439584;
ROM1[8568]<=26'd1948106; ROM2[8568]<=26'd11109866; ROM3[8568]<=26'd9699845; ROM4[8568]<=26'd23434592;
ROM1[8569]<=26'd1943741; ROM2[8569]<=26'd11110303; ROM3[8569]<=26'd9703897; ROM4[8569]<=26'd23435603;
ROM1[8570]<=26'd1944656; ROM2[8570]<=26'd11113734; ROM3[8570]<=26'd9709057; ROM4[8570]<=26'd23439798;
ROM1[8571]<=26'd1950945; ROM2[8571]<=26'd11117414; ROM3[8571]<=26'd9711028; ROM4[8571]<=26'd23441324;
ROM1[8572]<=26'd1959432; ROM2[8572]<=26'd11114834; ROM3[8572]<=26'd9705860; ROM4[8572]<=26'd23437933;
ROM1[8573]<=26'd1966376; ROM2[8573]<=26'd11112808; ROM3[8573]<=26'd9698330; ROM4[8573]<=26'd23435366;
ROM1[8574]<=26'd1961154; ROM2[8574]<=26'd11109415; ROM3[8574]<=26'd9697670; ROM4[8574]<=26'd23432442;
ROM1[8575]<=26'd1960289; ROM2[8575]<=26'd11117937; ROM3[8575]<=26'd9711262; ROM4[8575]<=26'd23441403;
ROM1[8576]<=26'd1958448; ROM2[8576]<=26'd11121805; ROM3[8576]<=26'd9719128; ROM4[8576]<=26'd23447563;
ROM1[8577]<=26'd1949513; ROM2[8577]<=26'd11114501; ROM3[8577]<=26'd9714468; ROM4[8577]<=26'd23441922;
ROM1[8578]<=26'd1940588; ROM2[8578]<=26'd11109940; ROM3[8578]<=26'd9712690; ROM4[8578]<=26'd23439002;
ROM1[8579]<=26'd1939247; ROM2[8579]<=26'd11106868; ROM3[8579]<=26'd9709288; ROM4[8579]<=26'd23436803;
ROM1[8580]<=26'd1944297; ROM2[8580]<=26'd11104788; ROM3[8580]<=26'd9702135; ROM4[8580]<=26'd23432795;
ROM1[8581]<=26'd1958793; ROM2[8581]<=26'd11109217; ROM3[8581]<=26'd9700700; ROM4[8581]<=26'd23436639;
ROM1[8582]<=26'd1964832; ROM2[8582]<=26'd11111520; ROM3[8582]<=26'd9702242; ROM4[8582]<=26'd23438947;
ROM1[8583]<=26'd1957352; ROM2[8583]<=26'd11109239; ROM3[8583]<=26'd9702669; ROM4[8583]<=26'd23436555;
ROM1[8584]<=26'd1949310; ROM2[8584]<=26'd11108022; ROM3[8584]<=26'd9704592; ROM4[8584]<=26'd23435647;
ROM1[8585]<=26'd1944882; ROM2[8585]<=26'd11107611; ROM3[8585]<=26'd9706034; ROM4[8585]<=26'd23435125;
ROM1[8586]<=26'd1939929; ROM2[8586]<=26'd11107897; ROM3[8586]<=26'd9706299; ROM4[8586]<=26'd23435307;
ROM1[8587]<=26'd1938753; ROM2[8587]<=26'd11107638; ROM3[8587]<=26'd9706537; ROM4[8587]<=26'd23435501;
ROM1[8588]<=26'd1948327; ROM2[8588]<=26'd11111307; ROM3[8588]<=26'd9707816; ROM4[8588]<=26'd23438131;
ROM1[8589]<=26'd1968064; ROM2[8589]<=26'd11120234; ROM3[8589]<=26'd9711641; ROM4[8589]<=26'd23443867;
ROM1[8590]<=26'd1979676; ROM2[8590]<=26'd11125700; ROM3[8590]<=26'd9716319; ROM4[8590]<=26'd23449128;
ROM1[8591]<=26'd1969481; ROM2[8591]<=26'd11117286; ROM3[8591]<=26'd9711183; ROM4[8591]<=26'd23441737;
ROM1[8592]<=26'd1960066; ROM2[8592]<=26'd11112545; ROM3[8592]<=26'd9712483; ROM4[8592]<=26'd23440966;
ROM1[8593]<=26'd1954251; ROM2[8593]<=26'd11111458; ROM3[8593]<=26'd9716432; ROM4[8593]<=26'd23443951;
ROM1[8594]<=26'd1945149; ROM2[8594]<=26'd11106566; ROM3[8594]<=26'd9714867; ROM4[8594]<=26'd23440048;
ROM1[8595]<=26'd1941812; ROM2[8595]<=26'd11105613; ROM3[8595]<=26'd9714709; ROM4[8595]<=26'd23439739;
ROM1[8596]<=26'd1946873; ROM2[8596]<=26'd11109624; ROM3[8596]<=26'd9715569; ROM4[8596]<=26'd23440960;
ROM1[8597]<=26'd1961062; ROM2[8597]<=26'd11115694; ROM3[8597]<=26'd9715379; ROM4[8597]<=26'd23443854;
ROM1[8598]<=26'd1969887; ROM2[8598]<=26'd11113186; ROM3[8598]<=26'd9705217; ROM4[8598]<=26'd23439179;
ROM1[8599]<=26'd1965815; ROM2[8599]<=26'd11108758; ROM3[8599]<=26'd9700462; ROM4[8599]<=26'd23435461;
ROM1[8600]<=26'd1960106; ROM2[8600]<=26'd11107964; ROM3[8600]<=26'd9701654; ROM4[8600]<=26'd23435765;
ROM1[8601]<=26'd1954706; ROM2[8601]<=26'd11108167; ROM3[8601]<=26'd9703665; ROM4[8601]<=26'd23435722;
ROM1[8602]<=26'd1955241; ROM2[8602]<=26'd11114003; ROM3[8602]<=26'd9709377; ROM4[8602]<=26'd23442408;
ROM1[8603]<=26'd1956228; ROM2[8603]<=26'd11119104; ROM3[8603]<=26'd9714666; ROM4[8603]<=26'd23446711;
ROM1[8604]<=26'd1956201; ROM2[8604]<=26'd11116300; ROM3[8604]<=26'd9713290; ROM4[8604]<=26'd23444779;
ROM1[8605]<=26'd1963271; ROM2[8605]<=26'd11112845; ROM3[8605]<=26'd9708015; ROM4[8605]<=26'd23443218;
ROM1[8606]<=26'd1978555; ROM2[8606]<=26'd11115624; ROM3[8606]<=26'd9704609; ROM4[8606]<=26'd23445027;
ROM1[8607]<=26'd1989681; ROM2[8607]<=26'd11121980; ROM3[8607]<=26'd9711809; ROM4[8607]<=26'd23453815;
ROM1[8608]<=26'd1988816; ROM2[8608]<=26'd11124756; ROM3[8608]<=26'd9718287; ROM4[8608]<=26'd23458999;
ROM1[8609]<=26'd1972914; ROM2[8609]<=26'd11117032; ROM3[8609]<=26'd9715660; ROM4[8609]<=26'd23452520;
ROM1[8610]<=26'd1967320; ROM2[8610]<=26'd11114840; ROM3[8610]<=26'd9718532; ROM4[8610]<=26'd23453513;
ROM1[8611]<=26'd1964906; ROM2[8611]<=26'd11117740; ROM3[8611]<=26'd9722125; ROM4[8611]<=26'd23456162;
ROM1[8612]<=26'd1957470; ROM2[8612]<=26'd11112809; ROM3[8612]<=26'd9715078; ROM4[8612]<=26'd23450400;
ROM1[8613]<=26'd1961987; ROM2[8613]<=26'd11111117; ROM3[8613]<=26'd9706287; ROM4[8613]<=26'd23448044;
ROM1[8614]<=26'd1973907; ROM2[8614]<=26'd11111268; ROM3[8614]<=26'd9700376; ROM4[8614]<=26'd23444853;
ROM1[8615]<=26'd1981326; ROM2[8615]<=26'd11113104; ROM3[8615]<=26'd9697983; ROM4[8615]<=26'd23445966;
ROM1[8616]<=26'd1977258; ROM2[8616]<=26'd11113936; ROM3[8616]<=26'd9698394; ROM4[8616]<=26'd23446752;
ROM1[8617]<=26'd1969056; ROM2[8617]<=26'd11112973; ROM3[8617]<=26'd9700536; ROM4[8617]<=26'd23445071;
ROM1[8618]<=26'd1961756; ROM2[8618]<=26'd11113082; ROM3[8618]<=26'd9702624; ROM4[8618]<=26'd23444176;
ROM1[8619]<=26'd1950122; ROM2[8619]<=26'd11106700; ROM3[8619]<=26'd9699257; ROM4[8619]<=26'd23438034;
ROM1[8620]<=26'd1944850; ROM2[8620]<=26'd11103774; ROM3[8620]<=26'd9700244; ROM4[8620]<=26'd23435968;
ROM1[8621]<=26'd1955239; ROM2[8621]<=26'd11109509; ROM3[8621]<=26'd9706887; ROM4[8621]<=26'd23440997;
ROM1[8622]<=26'd1966436; ROM2[8622]<=26'd11111240; ROM3[8622]<=26'd9704509; ROM4[8622]<=26'd23441121;
ROM1[8623]<=26'd1969269; ROM2[8623]<=26'd11106973; ROM3[8623]<=26'd9694672; ROM4[8623]<=26'd23436181;
ROM1[8624]<=26'd1969092; ROM2[8624]<=26'd11108570; ROM3[8624]<=26'd9696793; ROM4[8624]<=26'd23437389;
ROM1[8625]<=26'd1964283; ROM2[8625]<=26'd11110757; ROM3[8625]<=26'd9703405; ROM4[8625]<=26'd23439627;
ROM1[8626]<=26'd1955920; ROM2[8626]<=26'd11108790; ROM3[8626]<=26'd9707398; ROM4[8626]<=26'd23441285;
ROM1[8627]<=26'd1959952; ROM2[8627]<=26'd11118394; ROM3[8627]<=26'd9720291; ROM4[8627]<=26'd23452382;
ROM1[8628]<=26'd1969391; ROM2[8628]<=26'd11133012; ROM3[8628]<=26'd9734431; ROM4[8628]<=26'd23465316;
ROM1[8629]<=26'd1962204; ROM2[8629]<=26'd11125871; ROM3[8629]<=26'd9725426; ROM4[8629]<=26'd23457946;
ROM1[8630]<=26'd1957330; ROM2[8630]<=26'd11112347; ROM3[8630]<=26'd9708433; ROM4[8630]<=26'd23442013;
ROM1[8631]<=26'd1963534; ROM2[8631]<=26'd11107368; ROM3[8631]<=26'd9696415; ROM4[8631]<=26'd23434475;
ROM1[8632]<=26'd1961815; ROM2[8632]<=26'd11102899; ROM3[8632]<=26'd9690084; ROM4[8632]<=26'd23428898;
ROM1[8633]<=26'd1959223; ROM2[8633]<=26'd11105006; ROM3[8633]<=26'd9693938; ROM4[8633]<=26'd23430486;
ROM1[8634]<=26'd1958048; ROM2[8634]<=26'd11111618; ROM3[8634]<=26'd9703762; ROM4[8634]<=26'd23438818;
ROM1[8635]<=26'd1952878; ROM2[8635]<=26'd11108938; ROM3[8635]<=26'd9706683; ROM4[8635]<=26'd23437264;
ROM1[8636]<=26'd1939740; ROM2[8636]<=26'd11100606; ROM3[8636]<=26'd9703961; ROM4[8636]<=26'd23432140;
ROM1[8637]<=26'd1938011; ROM2[8637]<=26'd11099835; ROM3[8637]<=26'd9707835; ROM4[8637]<=26'd23434131;
ROM1[8638]<=26'd1949974; ROM2[8638]<=26'd11103714; ROM3[8638]<=26'd9711058; ROM4[8638]<=26'd23438059;
ROM1[8639]<=26'd1963691; ROM2[8639]<=26'd11103655; ROM3[8639]<=26'd9708884; ROM4[8639]<=26'd23438230;
ROM1[8640]<=26'd1969948; ROM2[8640]<=26'd11101299; ROM3[8640]<=26'd9707634; ROM4[8640]<=26'd23438083;
ROM1[8641]<=26'd1967948; ROM2[8641]<=26'd11102452; ROM3[8641]<=26'd9710765; ROM4[8641]<=26'd23440829;
ROM1[8642]<=26'd1959892; ROM2[8642]<=26'd11101221; ROM3[8642]<=26'd9713774; ROM4[8642]<=26'd23441427;
ROM1[8643]<=26'd1957300; ROM2[8643]<=26'd11103470; ROM3[8643]<=26'd9720926; ROM4[8643]<=26'd23444520;
ROM1[8644]<=26'd1955152; ROM2[8644]<=26'd11106482; ROM3[8644]<=26'd9724724; ROM4[8644]<=26'd23445520;
ROM1[8645]<=26'd1951899; ROM2[8645]<=26'd11106274; ROM3[8645]<=26'd9724144; ROM4[8645]<=26'd23444275;
ROM1[8646]<=26'd1961313; ROM2[8646]<=26'd11111757; ROM3[8646]<=26'd9725469; ROM4[8646]<=26'd23449664;
ROM1[8647]<=26'd1969026; ROM2[8647]<=26'd11110004; ROM3[8647]<=26'd9717287; ROM4[8647]<=26'd23446884;
ROM1[8648]<=26'd1975112; ROM2[8648]<=26'd11107748; ROM3[8648]<=26'd9708231; ROM4[8648]<=26'd23440876;
ROM1[8649]<=26'd1973618; ROM2[8649]<=26'd11107140; ROM3[8649]<=26'd9705997; ROM4[8649]<=26'd23440178;
ROM1[8650]<=26'd1968343; ROM2[8650]<=26'd11108934; ROM3[8650]<=26'd9709588; ROM4[8650]<=26'd23441986;
ROM1[8651]<=26'd1969555; ROM2[8651]<=26'd11118528; ROM3[8651]<=26'd9719442; ROM4[8651]<=26'd23449667;
ROM1[8652]<=26'd1962523; ROM2[8652]<=26'd11117969; ROM3[8652]<=26'd9719923; ROM4[8652]<=26'd23448957;
ROM1[8653]<=26'd1954385; ROM2[8653]<=26'd11115705; ROM3[8653]<=26'd9718311; ROM4[8653]<=26'd23445902;
ROM1[8654]<=26'd1953056; ROM2[8654]<=26'd11113868; ROM3[8654]<=26'd9716131; ROM4[8654]<=26'd23443678;
ROM1[8655]<=26'd1956748; ROM2[8655]<=26'd11109264; ROM3[8655]<=26'd9705083; ROM4[8655]<=26'd23435939;
ROM1[8656]<=26'd1969506; ROM2[8656]<=26'd11111164; ROM3[8656]<=26'd9699306; ROM4[8656]<=26'd23436781;
ROM1[8657]<=26'd1973549; ROM2[8657]<=26'd11112690; ROM3[8657]<=26'd9700797; ROM4[8657]<=26'd23439530;
ROM1[8658]<=26'd1964627; ROM2[8658]<=26'd11108836; ROM3[8658]<=26'd9699289; ROM4[8658]<=26'd23435670;
ROM1[8659]<=26'd1952052; ROM2[8659]<=26'd11103969; ROM3[8659]<=26'd9699364; ROM4[8659]<=26'd23433053;
ROM1[8660]<=26'd1949535; ROM2[8660]<=26'd11105405; ROM3[8660]<=26'd9705061; ROM4[8660]<=26'd23437056;
ROM1[8661]<=26'd1948543; ROM2[8661]<=26'd11110454; ROM3[8661]<=26'd9712406; ROM4[8661]<=26'd23441206;
ROM1[8662]<=26'd1947327; ROM2[8662]<=26'd11113776; ROM3[8662]<=26'd9714604; ROM4[8662]<=26'd23442326;
ROM1[8663]<=26'd1962647; ROM2[8663]<=26'd11123141; ROM3[8663]<=26'd9722131; ROM4[8663]<=26'd23453005;
ROM1[8664]<=26'd1983942; ROM2[8664]<=26'd11131227; ROM3[8664]<=26'd9727158; ROM4[8664]<=26'd23463105;
ROM1[8665]<=26'd1985301; ROM2[8665]<=26'd11124181; ROM3[8665]<=26'd9717064; ROM4[8665]<=26'd23457512;
ROM1[8666]<=26'd1970671; ROM2[8666]<=26'd11111290; ROM3[8666]<=26'd9707586; ROM4[8666]<=26'd23446213;
ROM1[8667]<=26'd1958043; ROM2[8667]<=26'd11105509; ROM3[8667]<=26'd9704946; ROM4[8667]<=26'd23440268;
ROM1[8668]<=26'd1949170; ROM2[8668]<=26'd11101923; ROM3[8668]<=26'd9705894; ROM4[8668]<=26'd23437270;
ROM1[8669]<=26'd1944686; ROM2[8669]<=26'd11102910; ROM3[8669]<=26'd9711155; ROM4[8669]<=26'd23439122;
ROM1[8670]<=26'd1944282; ROM2[8670]<=26'd11106370; ROM3[8670]<=26'd9716412; ROM4[8670]<=26'd23443934;
ROM1[8671]<=26'd1947848; ROM2[8671]<=26'd11105994; ROM3[8671]<=26'd9715374; ROM4[8671]<=26'd23444111;
ROM1[8672]<=26'd1958942; ROM2[8672]<=26'd11105597; ROM3[8672]<=26'd9709664; ROM4[8672]<=26'd23442074;
ROM1[8673]<=26'd1973423; ROM2[8673]<=26'd11109072; ROM3[8673]<=26'd9707624; ROM4[8673]<=26'd23445578;
ROM1[8674]<=26'd1978049; ROM2[8674]<=26'd11113621; ROM3[8674]<=26'd9712395; ROM4[8674]<=26'd23451910;
ROM1[8675]<=26'd1971545; ROM2[8675]<=26'd11112610; ROM3[8675]<=26'd9715130; ROM4[8675]<=26'd23452712;
ROM1[8676]<=26'd1960372; ROM2[8676]<=26'd11109459; ROM3[8676]<=26'd9713662; ROM4[8676]<=26'd23449424;
ROM1[8677]<=26'd1954634; ROM2[8677]<=26'd11109704; ROM3[8677]<=26'd9715052; ROM4[8677]<=26'd23449504;
ROM1[8678]<=26'd1952249; ROM2[8678]<=26'd11111745; ROM3[8678]<=26'd9718967; ROM4[8678]<=26'd23452306;
ROM1[8679]<=26'd1952650; ROM2[8679]<=26'd11110787; ROM3[8679]<=26'd9717147; ROM4[8679]<=26'd23452392;
ROM1[8680]<=26'd1960030; ROM2[8680]<=26'd11110273; ROM3[8680]<=26'd9711817; ROM4[8680]<=26'd23450789;
ROM1[8681]<=26'd1974474; ROM2[8681]<=26'd11112165; ROM3[8681]<=26'd9706676; ROM4[8681]<=26'd23450957;
ROM1[8682]<=26'd1979510; ROM2[8682]<=26'd11111349; ROM3[8682]<=26'd9705845; ROM4[8682]<=26'd23450171;
ROM1[8683]<=26'd1974346; ROM2[8683]<=26'd11111616; ROM3[8683]<=26'd9707753; ROM4[8683]<=26'd23450755;
ROM1[8684]<=26'd1968738; ROM2[8684]<=26'd11112118; ROM3[8684]<=26'd9712005; ROM4[8684]<=26'd23452212;
ROM1[8685]<=26'd1965191; ROM2[8685]<=26'd11113301; ROM3[8685]<=26'd9716879; ROM4[8685]<=26'd23453916;
ROM1[8686]<=26'd1964116; ROM2[8686]<=26'd11118768; ROM3[8686]<=26'd9724343; ROM4[8686]<=26'd23459598;
ROM1[8687]<=26'd1966058; ROM2[8687]<=26'd11122418; ROM3[8687]<=26'd9729277; ROM4[8687]<=26'd23462796;
ROM1[8688]<=26'd1968020; ROM2[8688]<=26'd11120331; ROM3[8688]<=26'd9723472; ROM4[8688]<=26'd23458841;
ROM1[8689]<=26'd1979216; ROM2[8689]<=26'd11120274; ROM3[8689]<=26'd9718152; ROM4[8689]<=26'd23456145;
ROM1[8690]<=26'd1985804; ROM2[8690]<=26'd11120236; ROM3[8690]<=26'd9714039; ROM4[8690]<=26'd23454760;
ROM1[8691]<=26'd1972747; ROM2[8691]<=26'd11110550; ROM3[8691]<=26'd9705403; ROM4[8691]<=26'd23445415;
ROM1[8692]<=26'd1964627; ROM2[8692]<=26'd11107557; ROM3[8692]<=26'd9707287; ROM4[8692]<=26'd23444269;
ROM1[8693]<=26'd1960820; ROM2[8693]<=26'd11107738; ROM3[8693]<=26'd9711716; ROM4[8693]<=26'd23446326;
ROM1[8694]<=26'd1952137; ROM2[8694]<=26'd11106710; ROM3[8694]<=26'd9712694; ROM4[8694]<=26'd23444949;
ROM1[8695]<=26'd1951469; ROM2[8695]<=26'd11109342; ROM3[8695]<=26'd9715741; ROM4[8695]<=26'd23445702;
ROM1[8696]<=26'd1958661; ROM2[8696]<=26'd11113277; ROM3[8696]<=26'd9718451; ROM4[8696]<=26'd23448893;
ROM1[8697]<=26'd1973070; ROM2[8697]<=26'd11120130; ROM3[8697]<=26'd9719593; ROM4[8697]<=26'd23452341;
ROM1[8698]<=26'd1988004; ROM2[8698]<=26'd11125439; ROM3[8698]<=26'd9719716; ROM4[8698]<=26'd23455692;
ROM1[8699]<=26'd1992942; ROM2[8699]<=26'd11130856; ROM3[8699]<=26'd9725673; ROM4[8699]<=26'd23463208;
ROM1[8700]<=26'd1986312; ROM2[8700]<=26'd11130308; ROM3[8700]<=26'd9729060; ROM4[8700]<=26'd23463758;
ROM1[8701]<=26'd1966395; ROM2[8701]<=26'd11117974; ROM3[8701]<=26'd9721478; ROM4[8701]<=26'd23452776;
ROM1[8702]<=26'd1951251; ROM2[8702]<=26'd11106661; ROM3[8702]<=26'd9714072; ROM4[8702]<=26'd23443427;
ROM1[8703]<=26'd1946517; ROM2[8703]<=26'd11105932; ROM3[8703]<=26'd9715317; ROM4[8703]<=26'd23442770;
ROM1[8704]<=26'd1948402; ROM2[8704]<=26'd11107073; ROM3[8704]<=26'd9714527; ROM4[8704]<=26'd23442810;
ROM1[8705]<=26'd1960929; ROM2[8705]<=26'd11110765; ROM3[8705]<=26'd9711486; ROM4[8705]<=26'd23445402;
ROM1[8706]<=26'd1975331; ROM2[8706]<=26'd11113369; ROM3[8706]<=26'd9708028; ROM4[8706]<=26'd23447194;
ROM1[8707]<=26'd1977494; ROM2[8707]<=26'd11114498; ROM3[8707]<=26'd9708136; ROM4[8707]<=26'd23448270;
ROM1[8708]<=26'd1975463; ROM2[8708]<=26'd11117974; ROM3[8708]<=26'd9713983; ROM4[8708]<=26'd23450595;
ROM1[8709]<=26'd1964249; ROM2[8709]<=26'd11112676; ROM3[8709]<=26'd9714507; ROM4[8709]<=26'd23446365;
ROM1[8710]<=26'd1953340; ROM2[8710]<=26'd11106750; ROM3[8710]<=26'd9710498; ROM4[8710]<=26'd23441954;
ROM1[8711]<=26'd1946453; ROM2[8711]<=26'd11104585; ROM3[8711]<=26'd9710081; ROM4[8711]<=26'd23439503;
ROM1[8712]<=26'd1944337; ROM2[8712]<=26'd11104289; ROM3[8712]<=26'd9710703; ROM4[8712]<=26'd23440082;
ROM1[8713]<=26'd1955009; ROM2[8713]<=26'd11108914; ROM3[8713]<=26'd9710977; ROM4[8713]<=26'd23445076;
ROM1[8714]<=26'd1970245; ROM2[8714]<=26'd11113011; ROM3[8714]<=26'd9708338; ROM4[8714]<=26'd23446245;
ROM1[8715]<=26'd1974001; ROM2[8715]<=26'd11111424; ROM3[8715]<=26'd9701500; ROM4[8715]<=26'd23442689;
ROM1[8716]<=26'd1964569; ROM2[8716]<=26'd11107123; ROM3[8716]<=26'd9694497; ROM4[8716]<=26'd23437480;
ROM1[8717]<=26'd1957216; ROM2[8717]<=26'd11107322; ROM3[8717]<=26'd9695740; ROM4[8717]<=26'd23437290;
ROM1[8718]<=26'd1952929; ROM2[8718]<=26'd11109994; ROM3[8718]<=26'd9700112; ROM4[8718]<=26'd23439888;
ROM1[8719]<=26'd1950443; ROM2[8719]<=26'd11111386; ROM3[8719]<=26'd9704430; ROM4[8719]<=26'd23442864;
ROM1[8720]<=26'd1948727; ROM2[8720]<=26'd11113024; ROM3[8720]<=26'd9707996; ROM4[8720]<=26'd23444651;
ROM1[8721]<=26'd1951083; ROM2[8721]<=26'd11113487; ROM3[8721]<=26'd9706310; ROM4[8721]<=26'd23443948;
ROM1[8722]<=26'd1965639; ROM2[8722]<=26'd11117676; ROM3[8722]<=26'd9704339; ROM4[8722]<=26'd23445410;
ROM1[8723]<=26'd1977669; ROM2[8723]<=26'd11121677; ROM3[8723]<=26'd9702548; ROM4[8723]<=26'd23446931;
ROM1[8724]<=26'd1974767; ROM2[8724]<=26'd11117920; ROM3[8724]<=26'd9699956; ROM4[8724]<=26'd23443961;
ROM1[8725]<=26'd1970828; ROM2[8725]<=26'd11117828; ROM3[8725]<=26'd9706249; ROM4[8725]<=26'd23445833;
ROM1[8726]<=26'd1969285; ROM2[8726]<=26'd11122373; ROM3[8726]<=26'd9716992; ROM4[8726]<=26'd23451020;
ROM1[8727]<=26'd1966218; ROM2[8727]<=26'd11123502; ROM3[8727]<=26'd9721396; ROM4[8727]<=26'd23453600;
ROM1[8728]<=26'd1963267; ROM2[8728]<=26'd11123666; ROM3[8728]<=26'd9726299; ROM4[8728]<=26'd23456489;
ROM1[8729]<=26'd1965619; ROM2[8729]<=26'd11124853; ROM3[8729]<=26'd9728600; ROM4[8729]<=26'd23457856;
ROM1[8730]<=26'd1971546; ROM2[8730]<=26'd11121781; ROM3[8730]<=26'd9723710; ROM4[8730]<=26'd23454816;
ROM1[8731]<=26'd1984406; ROM2[8731]<=26'd11123610; ROM3[8731]<=26'd9721646; ROM4[8731]<=26'd23455798;
ROM1[8732]<=26'd1999001; ROM2[8732]<=26'd11134789; ROM3[8732]<=26'd9732424; ROM4[8732]<=26'd23468717;
ROM1[8733]<=26'd1995133; ROM2[8733]<=26'd11136503; ROM3[8733]<=26'd9735655; ROM4[8733]<=26'd23470851;
ROM1[8734]<=26'd1977851; ROM2[8734]<=26'd11125110; ROM3[8734]<=26'd9729694; ROM4[8734]<=26'd23461443;
ROM1[8735]<=26'd1975501; ROM2[8735]<=26'd11125608; ROM3[8735]<=26'd9735336; ROM4[8735]<=26'd23463709;
ROM1[8736]<=26'd1967612; ROM2[8736]<=26'd11124153; ROM3[8736]<=26'd9737423; ROM4[8736]<=26'd23461398;
ROM1[8737]<=26'd1963098; ROM2[8737]<=26'd11118838; ROM3[8737]<=26'd9735167; ROM4[8737]<=26'd23457624;
ROM1[8738]<=26'd1975415; ROM2[8738]<=26'd11126378; ROM3[8738]<=26'd9738002; ROM4[8738]<=26'd23462766;
ROM1[8739]<=26'd1986008; ROM2[8739]<=26'd11127514; ROM3[8739]<=26'd9730806; ROM4[8739]<=26'd23460639;
ROM1[8740]<=26'd1989749; ROM2[8740]<=26'd11125115; ROM3[8740]<=26'd9722134; ROM4[8740]<=26'd23457243;
ROM1[8741]<=26'd1988197; ROM2[8741]<=26'd11127462; ROM3[8741]<=26'd9723657; ROM4[8741]<=26'd23459496;
ROM1[8742]<=26'd1982946; ROM2[8742]<=26'd11126813; ROM3[8742]<=26'd9727409; ROM4[8742]<=26'd23460973;
ROM1[8743]<=26'd1976315; ROM2[8743]<=26'd11124353; ROM3[8743]<=26'd9728619; ROM4[8743]<=26'd23460377;
ROM1[8744]<=26'd1971340; ROM2[8744]<=26'd11124412; ROM3[8744]<=26'd9730382; ROM4[8744]<=26'd23460970;
ROM1[8745]<=26'd1971433; ROM2[8745]<=26'd11127699; ROM3[8745]<=26'd9735314; ROM4[8745]<=26'd23463509;
ROM1[8746]<=26'd1974988; ROM2[8746]<=26'd11129817; ROM3[8746]<=26'd9732827; ROM4[8746]<=26'd23464035;
ROM1[8747]<=26'd1990375; ROM2[8747]<=26'd11135075; ROM3[8747]<=26'd9732340; ROM4[8747]<=26'd23465677;
ROM1[8748]<=26'd1997209; ROM2[8748]<=26'd11133485; ROM3[8748]<=26'd9724776; ROM4[8748]<=26'd23461043;
ROM1[8749]<=26'd1982615; ROM2[8749]<=26'd11123229; ROM3[8749]<=26'd9710778; ROM4[8749]<=26'd23448286;
ROM1[8750]<=26'd1971271; ROM2[8750]<=26'd11117220; ROM3[8750]<=26'd9708737; ROM4[8750]<=26'd23442113;
ROM1[8751]<=26'd1959746; ROM2[8751]<=26'd11113178; ROM3[8751]<=26'd9706114; ROM4[8751]<=26'd23436773;
ROM1[8752]<=26'd1953283; ROM2[8752]<=26'd11112163; ROM3[8752]<=26'd9706140; ROM4[8752]<=26'd23436374;
ROM1[8753]<=26'd1952728; ROM2[8753]<=26'd11114583; ROM3[8753]<=26'd9711474; ROM4[8753]<=26'd23439845;
ROM1[8754]<=26'd1953128; ROM2[8754]<=26'd11116868; ROM3[8754]<=26'd9709801; ROM4[8754]<=26'd23441614;
ROM1[8755]<=26'd1958647; ROM2[8755]<=26'd11115557; ROM3[8755]<=26'd9702633; ROM4[8755]<=26'd23439617;
ROM1[8756]<=26'd1970783; ROM2[8756]<=26'd11115942; ROM3[8756]<=26'd9696568; ROM4[8756]<=26'd23435907;
ROM1[8757]<=26'd1974965; ROM2[8757]<=26'd11118767; ROM3[8757]<=26'd9696187; ROM4[8757]<=26'd23436575;
ROM1[8758]<=26'd1969612; ROM2[8758]<=26'd11120452; ROM3[8758]<=26'd9700573; ROM4[8758]<=26'd23437397;
ROM1[8759]<=26'd1961258; ROM2[8759]<=26'd11119073; ROM3[8759]<=26'd9704740; ROM4[8759]<=26'd23437109;
ROM1[8760]<=26'd1956308; ROM2[8760]<=26'd11117091; ROM3[8760]<=26'd9707299; ROM4[8760]<=26'd23436426;
ROM1[8761]<=26'd1950994; ROM2[8761]<=26'd11115440; ROM3[8761]<=26'd9710302; ROM4[8761]<=26'd23435363;
ROM1[8762]<=26'd1953630; ROM2[8762]<=26'd11117069; ROM3[8762]<=26'd9713813; ROM4[8762]<=26'd23437485;
ROM1[8763]<=26'd1964488; ROM2[8763]<=26'd11122506; ROM3[8763]<=26'd9716498; ROM4[8763]<=26'd23443440;
ROM1[8764]<=26'd1971198; ROM2[8764]<=26'd11120126; ROM3[8764]<=26'd9709840; ROM4[8764]<=26'd23441485;
ROM1[8765]<=26'd1971303; ROM2[8765]<=26'd11112636; ROM3[8765]<=26'd9701183; ROM4[8765]<=26'd23435828;
ROM1[8766]<=26'd1965967; ROM2[8766]<=26'd11110758; ROM3[8766]<=26'd9700613; ROM4[8766]<=26'd23434990;
ROM1[8767]<=26'd1954324; ROM2[8767]<=26'd11106617; ROM3[8767]<=26'd9701400; ROM4[8767]<=26'd23432306;
ROM1[8768]<=26'd1948621; ROM2[8768]<=26'd11106036; ROM3[8768]<=26'd9705848; ROM4[8768]<=26'd23435108;
ROM1[8769]<=26'd1946939; ROM2[8769]<=26'd11109629; ROM3[8769]<=26'd9713494; ROM4[8769]<=26'd23440528;
ROM1[8770]<=26'd1946205; ROM2[8770]<=26'd11111833; ROM3[8770]<=26'd9719629; ROM4[8770]<=26'd23443525;
ROM1[8771]<=26'd1951103; ROM2[8771]<=26'd11112224; ROM3[8771]<=26'd9719353; ROM4[8771]<=26'd23443395;
ROM1[8772]<=26'd1959124; ROM2[8772]<=26'd11110709; ROM3[8772]<=26'd9709799; ROM4[8772]<=26'd23439543;
ROM1[8773]<=26'd1969342; ROM2[8773]<=26'd11114403; ROM3[8773]<=26'd9704736; ROM4[8773]<=26'd23439800;
ROM1[8774]<=26'd1974133; ROM2[8774]<=26'd11119723; ROM3[8774]<=26'd9711036; ROM4[8774]<=26'd23445053;
ROM1[8775]<=26'd1966492; ROM2[8775]<=26'd11115910; ROM3[8775]<=26'd9709942; ROM4[8775]<=26'd23442454;
ROM1[8776]<=26'd1957676; ROM2[8776]<=26'd11110708; ROM3[8776]<=26'd9710087; ROM4[8776]<=26'd23439343;
ROM1[8777]<=26'd1956120; ROM2[8777]<=26'd11113379; ROM3[8777]<=26'd9717416; ROM4[8777]<=26'd23445692;
ROM1[8778]<=26'd1951825; ROM2[8778]<=26'd11113920; ROM3[8778]<=26'd9717362; ROM4[8778]<=26'd23445152;
ROM1[8779]<=26'd1952553; ROM2[8779]<=26'd11113025; ROM3[8779]<=26'd9713974; ROM4[8779]<=26'd23442339;
ROM1[8780]<=26'd1964188; ROM2[8780]<=26'd11116931; ROM3[8780]<=26'd9712966; ROM4[8780]<=26'd23443952;
ROM1[8781]<=26'd1977980; ROM2[8781]<=26'd11118971; ROM3[8781]<=26'd9710209; ROM4[8781]<=26'd23445180;
ROM1[8782]<=26'd1978963; ROM2[8782]<=26'd11117159; ROM3[8782]<=26'd9708237; ROM4[8782]<=26'd23444940;
ROM1[8783]<=26'd1973129; ROM2[8783]<=26'd11119161; ROM3[8783]<=26'd9712658; ROM4[8783]<=26'd23447087;
ROM1[8784]<=26'd1977675; ROM2[8784]<=26'd11129882; ROM3[8784]<=26'd9727596; ROM4[8784]<=26'd23457846;
ROM1[8785]<=26'd1982603; ROM2[8785]<=26'd11137861; ROM3[8785]<=26'd9738059; ROM4[8785]<=26'd23466368;
ROM1[8786]<=26'd1964748; ROM2[8786]<=26'd11125614; ROM3[8786]<=26'd9730093; ROM4[8786]<=26'd23455035;
ROM1[8787]<=26'd1956821; ROM2[8787]<=26'd11116677; ROM3[8787]<=26'd9724816; ROM4[8787]<=26'd23449581;
ROM1[8788]<=26'd1961823; ROM2[8788]<=26'd11116636; ROM3[8788]<=26'd9722966; ROM4[8788]<=26'd23451008;
ROM1[8789]<=26'd1974526; ROM2[8789]<=26'd11118322; ROM3[8789]<=26'd9720491; ROM4[8789]<=26'd23452090;
ROM1[8790]<=26'd1991524; ROM2[8790]<=26'd11128618; ROM3[8790]<=26'd9728143; ROM4[8790]<=26'd23462914;
ROM1[8791]<=26'd1990697; ROM2[8791]<=26'd11133230; ROM3[8791]<=26'd9734916; ROM4[8791]<=26'd23467459;
ROM1[8792]<=26'd1980157; ROM2[8792]<=26'd11130516; ROM3[8792]<=26'd9736275; ROM4[8792]<=26'd23465997;
ROM1[8793]<=26'd1969296; ROM2[8793]<=26'd11124591; ROM3[8793]<=26'd9735031; ROM4[8793]<=26'd23462690;
ROM1[8794]<=26'd1958746; ROM2[8794]<=26'd11119256; ROM3[8794]<=26'd9734196; ROM4[8794]<=26'd23459362;
ROM1[8795]<=26'd1955413; ROM2[8795]<=26'd11118447; ROM3[8795]<=26'd9736325; ROM4[8795]<=26'd23459417;
ROM1[8796]<=26'd1960505; ROM2[8796]<=26'd11118958; ROM3[8796]<=26'd9737040; ROM4[8796]<=26'd23460003;
ROM1[8797]<=26'd1972183; ROM2[8797]<=26'd11121901; ROM3[8797]<=26'd9731487; ROM4[8797]<=26'd23460125;
ROM1[8798]<=26'd1984261; ROM2[8798]<=26'd11124102; ROM3[8798]<=26'd9726783; ROM4[8798]<=26'd23460061;
ROM1[8799]<=26'd1987066; ROM2[8799]<=26'd11126261; ROM3[8799]<=26'd9728323; ROM4[8799]<=26'd23461096;
ROM1[8800]<=26'd1983977; ROM2[8800]<=26'd11129715; ROM3[8800]<=26'd9731695; ROM4[8800]<=26'd23463127;
ROM1[8801]<=26'd1971711; ROM2[8801]<=26'd11122994; ROM3[8801]<=26'd9728799; ROM4[8801]<=26'd23457667;
ROM1[8802]<=26'd1962346; ROM2[8802]<=26'd11117946; ROM3[8802]<=26'd9725316; ROM4[8802]<=26'd23452004;
ROM1[8803]<=26'd1959698; ROM2[8803]<=26'd11120246; ROM3[8803]<=26'd9728902; ROM4[8803]<=26'd23454386;
ROM1[8804]<=26'd1958827; ROM2[8804]<=26'd11115925; ROM3[8804]<=26'd9725978; ROM4[8804]<=26'd23450803;
ROM1[8805]<=26'd1966465; ROM2[8805]<=26'd11114158; ROM3[8805]<=26'd9721814; ROM4[8805]<=26'd23447466;
ROM1[8806]<=26'd1982640; ROM2[8806]<=26'd11118163; ROM3[8806]<=26'd9721312; ROM4[8806]<=26'd23451861;
ROM1[8807]<=26'd1984334; ROM2[8807]<=26'd11117926; ROM3[8807]<=26'd9720443; ROM4[8807]<=26'd23453064;
ROM1[8808]<=26'd1979412; ROM2[8808]<=26'd11118221; ROM3[8808]<=26'd9724394; ROM4[8808]<=26'd23455979;
ROM1[8809]<=26'd1975714; ROM2[8809]<=26'd11120955; ROM3[8809]<=26'd9732583; ROM4[8809]<=26'd23459069;
ROM1[8810]<=26'd1971370; ROM2[8810]<=26'd11121863; ROM3[8810]<=26'd9737664; ROM4[8810]<=26'd23461310;
ROM1[8811]<=26'd1963580; ROM2[8811]<=26'd11117952; ROM3[8811]<=26'd9739620; ROM4[8811]<=26'd23461891;
ROM1[8812]<=26'd1963994; ROM2[8812]<=26'd11119400; ROM3[8812]<=26'd9742517; ROM4[8812]<=26'd23464874;
ROM1[8813]<=26'd1974565; ROM2[8813]<=26'd11124429; ROM3[8813]<=26'd9743031; ROM4[8813]<=26'd23468819;
ROM1[8814]<=26'd1988027; ROM2[8814]<=26'd11126025; ROM3[8814]<=26'd9738988; ROM4[8814]<=26'd23470318;
ROM1[8815]<=26'd1997611; ROM2[8815]<=26'd11130678; ROM3[8815]<=26'd9738509; ROM4[8815]<=26'd23472931;
ROM1[8816]<=26'd1986851; ROM2[8816]<=26'd11125542; ROM3[8816]<=26'd9735655; ROM4[8816]<=26'd23467330;
ROM1[8817]<=26'd1974304; ROM2[8817]<=26'd11119384; ROM3[8817]<=26'd9732760; ROM4[8817]<=26'd23462477;
ROM1[8818]<=26'd1965860; ROM2[8818]<=26'd11118964; ROM3[8818]<=26'd9731826; ROM4[8818]<=26'd23459800;
ROM1[8819]<=26'd1953239; ROM2[8819]<=26'd11111961; ROM3[8819]<=26'd9726314; ROM4[8819]<=26'd23451218;
ROM1[8820]<=26'd1950299; ROM2[8820]<=26'd11112402; ROM3[8820]<=26'd9723965; ROM4[8820]<=26'd23449211;
ROM1[8821]<=26'd1954262; ROM2[8821]<=26'd11113674; ROM3[8821]<=26'd9721214; ROM4[8821]<=26'd23448250;
ROM1[8822]<=26'd1963670; ROM2[8822]<=26'd11111559; ROM3[8822]<=26'd9715314; ROM4[8822]<=26'd23444981;
ROM1[8823]<=26'd1972866; ROM2[8823]<=26'd11113080; ROM3[8823]<=26'd9708043; ROM4[8823]<=26'd23444030;
ROM1[8824]<=26'd1969281; ROM2[8824]<=26'd11111343; ROM3[8824]<=26'd9703967; ROM4[8824]<=26'd23439768;
ROM1[8825]<=26'd1962814; ROM2[8825]<=26'd11110439; ROM3[8825]<=26'd9705569; ROM4[8825]<=26'd23439494;
ROM1[8826]<=26'd1957815; ROM2[8826]<=26'd11112001; ROM3[8826]<=26'd9709186; ROM4[8826]<=26'd23440386;
ROM1[8827]<=26'd1955779; ROM2[8827]<=26'd11114640; ROM3[8827]<=26'd9713804; ROM4[8827]<=26'd23444047;
ROM1[8828]<=26'd1954362; ROM2[8828]<=26'd11117212; ROM3[8828]<=26'd9718011; ROM4[8828]<=26'd23447980;
ROM1[8829]<=26'd1957409; ROM2[8829]<=26'd11121577; ROM3[8829]<=26'd9722245; ROM4[8829]<=26'd23450651;
ROM1[8830]<=26'd1964511; ROM2[8830]<=26'd11120034; ROM3[8830]<=26'd9717477; ROM4[8830]<=26'd23447856;
ROM1[8831]<=26'd1971108; ROM2[8831]<=26'd11113726; ROM3[8831]<=26'd9707196; ROM4[8831]<=26'd23442471;
ROM1[8832]<=26'd1971524; ROM2[8832]<=26'd11113659; ROM3[8832]<=26'd9706956; ROM4[8832]<=26'd23442996;
ROM1[8833]<=26'd1965444; ROM2[8833]<=26'd11113008; ROM3[8833]<=26'd9707887; ROM4[8833]<=26'd23443199;
ROM1[8834]<=26'd1954520; ROM2[8834]<=26'd11106797; ROM3[8834]<=26'd9705617; ROM4[8834]<=26'd23439657;
ROM1[8835]<=26'd1950546; ROM2[8835]<=26'd11108794; ROM3[8835]<=26'd9712624; ROM4[8835]<=26'd23440092;
ROM1[8836]<=26'd1948079; ROM2[8836]<=26'd11111774; ROM3[8836]<=26'd9720685; ROM4[8836]<=26'd23443109;
ROM1[8837]<=26'd1944091; ROM2[8837]<=26'd11108540; ROM3[8837]<=26'd9720309; ROM4[8837]<=26'd23442482;
ROM1[8838]<=26'd1953864; ROM2[8838]<=26'd11112869; ROM3[8838]<=26'd9723460; ROM4[8838]<=26'd23448089;
ROM1[8839]<=26'd1970864; ROM2[8839]<=26'd11117924; ROM3[8839]<=26'd9721546; ROM4[8839]<=26'd23450538;
ROM1[8840]<=26'd1975863; ROM2[8840]<=26'd11115433; ROM3[8840]<=26'd9717105; ROM4[8840]<=26'd23447178;
ROM1[8841]<=26'd1975452; ROM2[8841]<=26'd11118211; ROM3[8841]<=26'd9724213; ROM4[8841]<=26'd23451324;
ROM1[8842]<=26'd1975685; ROM2[8842]<=26'd11126347; ROM3[8842]<=26'd9735814; ROM4[8842]<=26'd23460342;
ROM1[8843]<=26'd1967978; ROM2[8843]<=26'd11122337; ROM3[8843]<=26'd9737254; ROM4[8843]<=26'd23459195;
ROM1[8844]<=26'd1958888; ROM2[8844]<=26'd11119210; ROM3[8844]<=26'd9736352; ROM4[8844]<=26'd23457141;
ROM1[8845]<=26'd1955029; ROM2[8845]<=26'd11118263; ROM3[8845]<=26'd9734554; ROM4[8845]<=26'd23454945;
ROM1[8846]<=26'd1957648; ROM2[8846]<=26'd11116949; ROM3[8846]<=26'd9729904; ROM4[8846]<=26'd23451984;
ROM1[8847]<=26'd1969236; ROM2[8847]<=26'd11118829; ROM3[8847]<=26'd9725034; ROM4[8847]<=26'd23451291;
ROM1[8848]<=26'd1980222; ROM2[8848]<=26'd11121674; ROM3[8848]<=26'd9720013; ROM4[8848]<=26'd23451160;
ROM1[8849]<=26'd1979471; ROM2[8849]<=26'd11123187; ROM3[8849]<=26'd9720418; ROM4[8849]<=26'd23452525;
ROM1[8850]<=26'd1976218; ROM2[8850]<=26'd11127024; ROM3[8850]<=26'd9726621; ROM4[8850]<=26'd23457844;
ROM1[8851]<=26'd1975852; ROM2[8851]<=26'd11132206; ROM3[8851]<=26'd9735350; ROM4[8851]<=26'd23464378;
ROM1[8852]<=26'd1967596; ROM2[8852]<=26'd11126661; ROM3[8852]<=26'd9732683; ROM4[8852]<=26'd23461030;
ROM1[8853]<=26'd1958677; ROM2[8853]<=26'd11123864; ROM3[8853]<=26'd9729996; ROM4[8853]<=26'd23456674;
ROM1[8854]<=26'd1954910; ROM2[8854]<=26'd11119722; ROM3[8854]<=26'd9724939; ROM4[8854]<=26'd23450475;
ROM1[8855]<=26'd1959798; ROM2[8855]<=26'd11118968; ROM3[8855]<=26'd9718136; ROM4[8855]<=26'd23448469;
ROM1[8856]<=26'd1976087; ROM2[8856]<=26'd11125265; ROM3[8856]<=26'd9715376; ROM4[8856]<=26'd23452299;
ROM1[8857]<=26'd1979084; ROM2[8857]<=26'd11122868; ROM3[8857]<=26'd9709752; ROM4[8857]<=26'd23447811;
ROM1[8858]<=26'd1972242; ROM2[8858]<=26'd11120657; ROM3[8858]<=26'd9707733; ROM4[8858]<=26'd23444238;
ROM1[8859]<=26'd1968293; ROM2[8859]<=26'd11121902; ROM3[8859]<=26'd9713598; ROM4[8859]<=26'd23445257;
ROM1[8860]<=26'd1963125; ROM2[8860]<=26'd11119283; ROM3[8860]<=26'd9718281; ROM4[8860]<=26'd23445048;
ROM1[8861]<=26'd1953270; ROM2[8861]<=26'd11116043; ROM3[8861]<=26'd9721953; ROM4[8861]<=26'd23445076;
ROM1[8862]<=26'd1951178; ROM2[8862]<=26'd11115755; ROM3[8862]<=26'd9724191; ROM4[8862]<=26'd23447433;
ROM1[8863]<=26'd1956632; ROM2[8863]<=26'd11117083; ROM3[8863]<=26'd9718753; ROM4[8863]<=26'd23445645;
ROM1[8864]<=26'd1969146; ROM2[8864]<=26'd11118734; ROM3[8864]<=26'd9714480; ROM4[8864]<=26'd23444171;
ROM1[8865]<=26'd1975964; ROM2[8865]<=26'd11118705; ROM3[8865]<=26'd9710170; ROM4[8865]<=26'd23443545;
ROM1[8866]<=26'd1969677; ROM2[8866]<=26'd11117009; ROM3[8866]<=26'd9708292; ROM4[8866]<=26'd23440834;
ROM1[8867]<=26'd1964306; ROM2[8867]<=26'd11119124; ROM3[8867]<=26'd9716444; ROM4[8867]<=26'd23444845;
ROM1[8868]<=26'd1969066; ROM2[8868]<=26'd11128794; ROM3[8868]<=26'd9728845; ROM4[8868]<=26'd23455224;
ROM1[8869]<=26'd1963313; ROM2[8869]<=26'd11127979; ROM3[8869]<=26'd9730653; ROM4[8869]<=26'd23456182;
ROM1[8870]<=26'd1952407; ROM2[8870]<=26'd11119483; ROM3[8870]<=26'd9722334; ROM4[8870]<=26'd23447544;
ROM1[8871]<=26'd1950354; ROM2[8871]<=26'd11113121; ROM3[8871]<=26'd9713767; ROM4[8871]<=26'd23442384;
ROM1[8872]<=26'd1957209; ROM2[8872]<=26'd11112160; ROM3[8872]<=26'd9707148; ROM4[8872]<=26'd23439615;
ROM1[8873]<=26'd1968853; ROM2[8873]<=26'd11115445; ROM3[8873]<=26'd9703787; ROM4[8873]<=26'd23440547;
ROM1[8874]<=26'd1975639; ROM2[8874]<=26'd11120361; ROM3[8874]<=26'd9710494; ROM4[8874]<=26'd23446750;
ROM1[8875]<=26'd1973376; ROM2[8875]<=26'd11123484; ROM3[8875]<=26'd9716915; ROM4[8875]<=26'd23450179;
ROM1[8876]<=26'd1958895; ROM2[8876]<=26'd11115904; ROM3[8876]<=26'd9712436; ROM4[8876]<=26'd23443389;
ROM1[8877]<=26'd1952151; ROM2[8877]<=26'd11113546; ROM3[8877]<=26'd9714010; ROM4[8877]<=26'd23442457;
ROM1[8878]<=26'd1948248; ROM2[8878]<=26'd11114528; ROM3[8878]<=26'd9718374; ROM4[8878]<=26'd23443231;
ROM1[8879]<=26'd1948997; ROM2[8879]<=26'd11111247; ROM3[8879]<=26'd9714764; ROM4[8879]<=26'd23440072;
ROM1[8880]<=26'd1958982; ROM2[8880]<=26'd11109976; ROM3[8880]<=26'd9709230; ROM4[8880]<=26'd23439160;
ROM1[8881]<=26'd1971814; ROM2[8881]<=26'd11112623; ROM3[8881]<=26'd9706603; ROM4[8881]<=26'd23441151;
ROM1[8882]<=26'd1976290; ROM2[8882]<=26'd11116401; ROM3[8882]<=26'd9709142; ROM4[8882]<=26'd23443250;
ROM1[8883]<=26'd1969282; ROM2[8883]<=26'd11117685; ROM3[8883]<=26'd9711781; ROM4[8883]<=26'd23444080;
ROM1[8884]<=26'd1960537; ROM2[8884]<=26'd11115815; ROM3[8884]<=26'd9714836; ROM4[8884]<=26'd23443933;
ROM1[8885]<=26'd1959070; ROM2[8885]<=26'd11117550; ROM3[8885]<=26'd9718501; ROM4[8885]<=26'd23446543;
ROM1[8886]<=26'd1961932; ROM2[8886]<=26'd11125248; ROM3[8886]<=26'd9727665; ROM4[8886]<=26'd23454470;
ROM1[8887]<=26'd1960930; ROM2[8887]<=26'd11123741; ROM3[8887]<=26'd9726729; ROM4[8887]<=26'd23453261;
ROM1[8888]<=26'd1961915; ROM2[8888]<=26'd11118086; ROM3[8888]<=26'd9717123; ROM4[8888]<=26'd23446897;
ROM1[8889]<=26'd1972334; ROM2[8889]<=26'd11116644; ROM3[8889]<=26'd9709954; ROM4[8889]<=26'd23442920;
ROM1[8890]<=26'd1973340; ROM2[8890]<=26'd11111476; ROM3[8890]<=26'd9701451; ROM4[8890]<=26'd23437431;
ROM1[8891]<=26'd1968571; ROM2[8891]<=26'd11111321; ROM3[8891]<=26'd9701439; ROM4[8891]<=26'd23436884;
ROM1[8892]<=26'd1969451; ROM2[8892]<=26'd11119179; ROM3[8892]<=26'd9712180; ROM4[8892]<=26'd23445824;
ROM1[8893]<=26'd1970954; ROM2[8893]<=26'd11126926; ROM3[8893]<=26'd9722596; ROM4[8893]<=26'd23453773;
ROM1[8894]<=26'd1963913; ROM2[8894]<=26'd11124811; ROM3[8894]<=26'd9723885; ROM4[8894]<=26'd23453157;
ROM1[8895]<=26'd1962732; ROM2[8895]<=26'd11124883; ROM3[8895]<=26'd9727247; ROM4[8895]<=26'd23453947;
ROM1[8896]<=26'd1971280; ROM2[8896]<=26'd11131035; ROM3[8896]<=26'd9731020; ROM4[8896]<=26'd23458091;
ROM1[8897]<=26'd1976133; ROM2[8897]<=26'd11126410; ROM3[8897]<=26'd9720549; ROM4[8897]<=26'd23451768;
ROM1[8898]<=26'd1984999; ROM2[8898]<=26'd11124848; ROM3[8898]<=26'd9716138; ROM4[8898]<=26'd23451002;
ROM1[8899]<=26'd1983317; ROM2[8899]<=26'd11123782; ROM3[8899]<=26'd9717889; ROM4[8899]<=26'd23452376;
ROM1[8900]<=26'd1984493; ROM2[8900]<=26'd11129671; ROM3[8900]<=26'd9725652; ROM4[8900]<=26'd23457400;
ROM1[8901]<=26'd1986554; ROM2[8901]<=26'd11135066; ROM3[8901]<=26'd9734017; ROM4[8901]<=26'd23463486;
ROM1[8902]<=26'd1967935; ROM2[8902]<=26'd11121956; ROM3[8902]<=26'd9722828; ROM4[8902]<=26'd23451314;
ROM1[8903]<=26'd1957248; ROM2[8903]<=26'd11114276; ROM3[8903]<=26'd9719983; ROM4[8903]<=26'd23443835;
ROM1[8904]<=26'd1955463; ROM2[8904]<=26'd11110301; ROM3[8904]<=26'd9716270; ROM4[8904]<=26'd23439677;
ROM1[8905]<=26'd1962095; ROM2[8905]<=26'd11110286; ROM3[8905]<=26'd9711022; ROM4[8905]<=26'd23438353;
ROM1[8906]<=26'd1985989; ROM2[8906]<=26'd11123830; ROM3[8906]<=26'd9717522; ROM4[8906]<=26'd23449184;
ROM1[8907]<=26'd1991666; ROM2[8907]<=26'd11129337; ROM3[8907]<=26'd9717970; ROM4[8907]<=26'd23452442;
ROM1[8908]<=26'd1975389; ROM2[8908]<=26'd11120100; ROM3[8908]<=26'd9710485; ROM4[8908]<=26'd23443019;
ROM1[8909]<=26'd1964063; ROM2[8909]<=26'd11116542; ROM3[8909]<=26'd9709720; ROM4[8909]<=26'd23438744;
ROM1[8910]<=26'd1962160; ROM2[8910]<=26'd11119731; ROM3[8910]<=26'd9713459; ROM4[8910]<=26'd23441667;
ROM1[8911]<=26'd1956816; ROM2[8911]<=26'd11119760; ROM3[8911]<=26'd9715780; ROM4[8911]<=26'd23443322;
ROM1[8912]<=26'd1953716; ROM2[8912]<=26'd11117677; ROM3[8912]<=26'd9713419; ROM4[8912]<=26'd23441635;
ROM1[8913]<=26'd1956131; ROM2[8913]<=26'd11114025; ROM3[8913]<=26'd9706770; ROM4[8913]<=26'd23436720;
ROM1[8914]<=26'd1964852; ROM2[8914]<=26'd11112792; ROM3[8914]<=26'd9699041; ROM4[8914]<=26'd23433515;
ROM1[8915]<=26'd1973398; ROM2[8915]<=26'd11115636; ROM3[8915]<=26'd9696929; ROM4[8915]<=26'd23434274;
ROM1[8916]<=26'd1970005; ROM2[8916]<=26'd11116326; ROM3[8916]<=26'd9700644; ROM4[8916]<=26'd23437240;
ROM1[8917]<=26'd1958412; ROM2[8917]<=26'd11113112; ROM3[8917]<=26'd9700926; ROM4[8917]<=26'd23434947;
ROM1[8918]<=26'd1950872; ROM2[8918]<=26'd11110264; ROM3[8918]<=26'd9701700; ROM4[8918]<=26'd23431272;
ROM1[8919]<=26'd1942801; ROM2[8919]<=26'd11106849; ROM3[8919]<=26'd9701691; ROM4[8919]<=26'd23428523;
ROM1[8920]<=26'd1945395; ROM2[8920]<=26'd11110913; ROM3[8920]<=26'd9707234; ROM4[8920]<=26'd23431496;
ROM1[8921]<=26'd1955311; ROM2[8921]<=26'd11116046; ROM3[8921]<=26'd9710231; ROM4[8921]<=26'd23436721;
ROM1[8922]<=26'd1962446; ROM2[8922]<=26'd11113769; ROM3[8922]<=26'd9701900; ROM4[8922]<=26'd23432216;
ROM1[8923]<=26'd1966957; ROM2[8923]<=26'd11110278; ROM3[8923]<=26'd9692290; ROM4[8923]<=26'd23427357;
ROM1[8924]<=26'd1963945; ROM2[8924]<=26'd11109154; ROM3[8924]<=26'd9689348; ROM4[8924]<=26'd23426803;
ROM1[8925]<=26'd1957384; ROM2[8925]<=26'd11107915; ROM3[8925]<=26'd9692041; ROM4[8925]<=26'd23427117;
ROM1[8926]<=26'd1952238; ROM2[8926]<=26'd11108699; ROM3[8926]<=26'd9695636; ROM4[8926]<=26'd23427586;
ROM1[8927]<=26'd1950558; ROM2[8927]<=26'd11110452; ROM3[8927]<=26'd9699027; ROM4[8927]<=26'd23430418;
ROM1[8928]<=26'd1945971; ROM2[8928]<=26'd11108930; ROM3[8928]<=26'd9700429; ROM4[8928]<=26'd23431356;
ROM1[8929]<=26'd1946748; ROM2[8929]<=26'd11108730; ROM3[8929]<=26'd9700574; ROM4[8929]<=26'd23431272;
ROM1[8930]<=26'd1957282; ROM2[8930]<=26'd11109622; ROM3[8930]<=26'd9699410; ROM4[8930]<=26'd23432575;
ROM1[8931]<=26'd1972709; ROM2[8931]<=26'd11116065; ROM3[8931]<=26'd9698533; ROM4[8931]<=26'd23437213;
ROM1[8932]<=26'd1977888; ROM2[8932]<=26'd11121399; ROM3[8932]<=26'd9701584; ROM4[8932]<=26'd23441080;
ROM1[8933]<=26'd1979037; ROM2[8933]<=26'd11125709; ROM3[8933]<=26'd9709267; ROM4[8933]<=26'd23445590;
ROM1[8934]<=26'd1972670; ROM2[8934]<=26'd11124651; ROM3[8934]<=26'd9713514; ROM4[8934]<=26'd23448411;
ROM1[8935]<=26'd1964214; ROM2[8935]<=26'd11120914; ROM3[8935]<=26'd9715817; ROM4[8935]<=26'd23447250;
ROM1[8936]<=26'd1963965; ROM2[8936]<=26'd11125627; ROM3[8936]<=26'd9725057; ROM4[8936]<=26'd23452046;
ROM1[8937]<=26'd1961640; ROM2[8937]<=26'd11123646; ROM3[8937]<=26'd9725415; ROM4[8937]<=26'd23450568;
ROM1[8938]<=26'd1959677; ROM2[8938]<=26'd11115136; ROM3[8938]<=26'd9715552; ROM4[8938]<=26'd23441945;
ROM1[8939]<=26'd1973212; ROM2[8939]<=26'd11115223; ROM3[8939]<=26'd9708927; ROM4[8939]<=26'd23439941;
ROM1[8940]<=26'd1975410; ROM2[8940]<=26'd11110892; ROM3[8940]<=26'd9704161; ROM4[8940]<=26'd23436290;
ROM1[8941]<=26'd1966327; ROM2[8941]<=26'd11108150; ROM3[8941]<=26'd9702962; ROM4[8941]<=26'd23433765;
ROM1[8942]<=26'd1965882; ROM2[8942]<=26'd11114118; ROM3[8942]<=26'd9712013; ROM4[8942]<=26'd23440448;
ROM1[8943]<=26'd1960959; ROM2[8943]<=26'd11112505; ROM3[8943]<=26'd9716950; ROM4[8943]<=26'd23441952;
ROM1[8944]<=26'd1951216; ROM2[8944]<=26'd11109561; ROM3[8944]<=26'd9715239; ROM4[8944]<=26'd23439645;
ROM1[8945]<=26'd1951398; ROM2[8945]<=26'd11110835; ROM3[8945]<=26'd9716977; ROM4[8945]<=26'd23441155;
ROM1[8946]<=26'd1959733; ROM2[8946]<=26'd11115023; ROM3[8946]<=26'd9719043; ROM4[8946]<=26'd23444774;
ROM1[8947]<=26'd1971093; ROM2[8947]<=26'd11119496; ROM3[8947]<=26'd9716420; ROM4[8947]<=26'd23446499;
ROM1[8948]<=26'd1979173; ROM2[8948]<=26'd11119101; ROM3[8948]<=26'd9710063; ROM4[8948]<=26'd23444510;
ROM1[8949]<=26'd1977925; ROM2[8949]<=26'd11119318; ROM3[8949]<=26'd9711304; ROM4[8949]<=26'd23445189;
ROM1[8950]<=26'd1971345; ROM2[8950]<=26'd11119800; ROM3[8950]<=26'd9715225; ROM4[8950]<=26'd23445008;
ROM1[8951]<=26'd1965690; ROM2[8951]<=26'd11119967; ROM3[8951]<=26'd9719986; ROM4[8951]<=26'd23446362;
ROM1[8952]<=26'd1964031; ROM2[8952]<=26'd11122980; ROM3[8952]<=26'd9725374; ROM4[8952]<=26'd23451591;
ROM1[8953]<=26'd1969977; ROM2[8953]<=26'd11131477; ROM3[8953]<=26'd9737083; ROM4[8953]<=26'd23461747;
ROM1[8954]<=26'd1981014; ROM2[8954]<=26'd11140579; ROM3[8954]<=26'd9744209; ROM4[8954]<=26'd23470902;
ROM1[8955]<=26'd1981551; ROM2[8955]<=26'd11132775; ROM3[8955]<=26'd9729474; ROM4[8955]<=26'd23460975;
ROM1[8956]<=26'd1983401; ROM2[8956]<=26'd11121761; ROM3[8956]<=26'd9712914; ROM4[8956]<=26'd23447401;
ROM1[8957]<=26'd1980822; ROM2[8957]<=26'd11119385; ROM3[8957]<=26'd9708036; ROM4[8957]<=26'd23443599;
ROM1[8958]<=26'd1972880; ROM2[8958]<=26'd11118074; ROM3[8958]<=26'd9707051; ROM4[8958]<=26'd23441400;
ROM1[8959]<=26'd1969819; ROM2[8959]<=26'd11121608; ROM3[8959]<=26'd9714912; ROM4[8959]<=26'd23445768;
ROM1[8960]<=26'd1969887; ROM2[8960]<=26'd11126716; ROM3[8960]<=26'd9724002; ROM4[8960]<=26'd23452482;
ROM1[8961]<=26'd1959387; ROM2[8961]<=26'd11121728; ROM3[8961]<=26'd9722756; ROM4[8961]<=26'd23448974;
ROM1[8962]<=26'd1954086; ROM2[8962]<=26'd11118333; ROM3[8962]<=26'd9719151; ROM4[8962]<=26'd23446758;
ROM1[8963]<=26'd1965917; ROM2[8963]<=26'd11123488; ROM3[8963]<=26'd9719697; ROM4[8963]<=26'd23450379;
ROM1[8964]<=26'd1979335; ROM2[8964]<=26'd11123538; ROM3[8964]<=26'd9715333; ROM4[8964]<=26'd23449018;
ROM1[8965]<=26'd1984265; ROM2[8965]<=26'd11123539; ROM3[8965]<=26'd9710672; ROM4[8965]<=26'd23450001;
ROM1[8966]<=26'd1980670; ROM2[8966]<=26'd11125322; ROM3[8966]<=26'd9715409; ROM4[8966]<=26'd23452387;
ROM1[8967]<=26'd1974625; ROM2[8967]<=26'd11124673; ROM3[8967]<=26'd9721647; ROM4[8967]<=26'd23454824;
ROM1[8968]<=26'd1965417; ROM2[8968]<=26'd11120272; ROM3[8968]<=26'd9720973; ROM4[8968]<=26'd23451722;
ROM1[8969]<=26'd1957204; ROM2[8969]<=26'd11117748; ROM3[8969]<=26'd9721662; ROM4[8969]<=26'd23449104;
ROM1[8970]<=26'd1954293; ROM2[8970]<=26'd11117303; ROM3[8970]<=26'd9723970; ROM4[8970]<=26'd23450495;
ROM1[8971]<=26'd1951047; ROM2[8971]<=26'd11112331; ROM3[8971]<=26'd9717073; ROM4[8971]<=26'd23443498;
ROM1[8972]<=26'd1961138; ROM2[8972]<=26'd11113144; ROM3[8972]<=26'd9712223; ROM4[8972]<=26'd23442067;
ROM1[8973]<=26'd1972745; ROM2[8973]<=26'd11114553; ROM3[8973]<=26'd9707924; ROM4[8973]<=26'd23442370;
ROM1[8974]<=26'd1970705; ROM2[8974]<=26'd11113013; ROM3[8974]<=26'd9706613; ROM4[8974]<=26'd23440373;
ROM1[8975]<=26'd1967978; ROM2[8975]<=26'd11117037; ROM3[8975]<=26'd9714217; ROM4[8975]<=26'd23443731;
ROM1[8976]<=26'd1968380; ROM2[8976]<=26'd11123078; ROM3[8976]<=26'd9725216; ROM4[8976]<=26'd23450955;
ROM1[8977]<=26'd1966478; ROM2[8977]<=26'd11125695; ROM3[8977]<=26'd9730667; ROM4[8977]<=26'd23454848;
ROM1[8978]<=26'd1954316; ROM2[8978]<=26'd11117763; ROM3[8978]<=26'd9724029; ROM4[8978]<=26'd23446488;
ROM1[8979]<=26'd1954807; ROM2[8979]<=26'd11116824; ROM3[8979]<=26'd9721790; ROM4[8979]<=26'd23443975;
ROM1[8980]<=26'd1965153; ROM2[8980]<=26'd11120512; ROM3[8980]<=26'd9720178; ROM4[8980]<=26'd23445715;
ROM1[8981]<=26'd1973006; ROM2[8981]<=26'd11117860; ROM3[8981]<=26'd9711777; ROM4[8981]<=26'd23441088;
ROM1[8982]<=26'd1976784; ROM2[8982]<=26'd11119478; ROM3[8982]<=26'd9711804; ROM4[8982]<=26'd23441930;
ROM1[8983]<=26'd1975742; ROM2[8983]<=26'd11124571; ROM3[8983]<=26'd9719230; ROM4[8983]<=26'd23448360;
ROM1[8984]<=26'd1974852; ROM2[8984]<=26'd11129023; ROM3[8984]<=26'd9727138; ROM4[8984]<=26'd23453824;
ROM1[8985]<=26'd1965674; ROM2[8985]<=26'd11123878; ROM3[8985]<=26'd9725152; ROM4[8985]<=26'd23449232;
ROM1[8986]<=26'd1953205; ROM2[8986]<=26'd11117725; ROM3[8986]<=26'd9721230; ROM4[8986]<=26'd23444134;
ROM1[8987]<=26'd1949776; ROM2[8987]<=26'd11114737; ROM3[8987]<=26'd9718554; ROM4[8987]<=26'd23442357;
ROM1[8988]<=26'd1952021; ROM2[8988]<=26'd11113257; ROM3[8988]<=26'd9711786; ROM4[8988]<=26'd23438739;
ROM1[8989]<=26'd1965395; ROM2[8989]<=26'd11117051; ROM3[8989]<=26'd9707414; ROM4[8989]<=26'd23440310;
ROM1[8990]<=26'd1975833; ROM2[8990]<=26'd11119278; ROM3[8990]<=26'd9706159; ROM4[8990]<=26'd23442647;
ROM1[8991]<=26'd1974318; ROM2[8991]<=26'd11118565; ROM3[8991]<=26'd9706616; ROM4[8991]<=26'd23442992;
ROM1[8992]<=26'd1965402; ROM2[8992]<=26'd11115398; ROM3[8992]<=26'd9706843; ROM4[8992]<=26'd23441818;
ROM1[8993]<=26'd1964329; ROM2[8993]<=26'd11118633; ROM3[8993]<=26'd9714440; ROM4[8993]<=26'd23445726;
ROM1[8994]<=26'd1965210; ROM2[8994]<=26'd11124963; ROM3[8994]<=26'd9726354; ROM4[8994]<=26'd23454683;
ROM1[8995]<=26'd1963865; ROM2[8995]<=26'd11125985; ROM3[8995]<=26'd9730173; ROM4[8995]<=26'd23456805;
ROM1[8996]<=26'd1965391; ROM2[8996]<=26'd11122238; ROM3[8996]<=26'd9726977; ROM4[8996]<=26'd23453376;
ROM1[8997]<=26'd1972573; ROM2[8997]<=26'd11118456; ROM3[8997]<=26'd9718119; ROM4[8997]<=26'd23448859;
ROM1[8998]<=26'd1980599; ROM2[8998]<=26'd11117607; ROM3[8998]<=26'd9710785; ROM4[8998]<=26'd23445109;
ROM1[8999]<=26'd1982953; ROM2[8999]<=26'd11124108; ROM3[8999]<=26'd9716530; ROM4[8999]<=26'd23451075;
ROM1[9000]<=26'd1979990; ROM2[9000]<=26'd11128589; ROM3[9000]<=26'd9722380; ROM4[9000]<=26'd23456003;
ROM1[9001]<=26'd1966566; ROM2[9001]<=26'd11120821; ROM3[9001]<=26'd9717929; ROM4[9001]<=26'd23448673;
ROM1[9002]<=26'd1957112; ROM2[9002]<=26'd11118287; ROM3[9002]<=26'd9717634; ROM4[9002]<=26'd23445789;
ROM1[9003]<=26'd1954832; ROM2[9003]<=26'd11121150; ROM3[9003]<=26'd9721126; ROM4[9003]<=26'd23448809;
ROM1[9004]<=26'd1959159; ROM2[9004]<=26'd11124468; ROM3[9004]<=26'd9721550; ROM4[9004]<=26'd23449439;
ROM1[9005]<=26'd1967000; ROM2[9005]<=26'd11123751; ROM3[9005]<=26'd9717203; ROM4[9005]<=26'd23446829;
ROM1[9006]<=26'd1977047; ROM2[9006]<=26'd11122869; ROM3[9006]<=26'd9710965; ROM4[9006]<=26'd23445358;
ROM1[9007]<=26'd1975666; ROM2[9007]<=26'd11118965; ROM3[9007]<=26'd9705177; ROM4[9007]<=26'd23440720;
ROM1[9008]<=26'd1968382; ROM2[9008]<=26'd11114699; ROM3[9008]<=26'd9705987; ROM4[9008]<=26'd23438546;
ROM1[9009]<=26'd1967286; ROM2[9009]<=26'd11120362; ROM3[9009]<=26'd9717928; ROM4[9009]<=26'd23446815;
ROM1[9010]<=26'd1966096; ROM2[9010]<=26'd11122917; ROM3[9010]<=26'd9724137; ROM4[9010]<=26'd23451077;
ROM1[9011]<=26'd1956027; ROM2[9011]<=26'd11119212; ROM3[9011]<=26'd9725437; ROM4[9011]<=26'd23447629;
ROM1[9012]<=26'd1950966; ROM2[9012]<=26'd11117268; ROM3[9012]<=26'd9725035; ROM4[9012]<=26'd23444569;
ROM1[9013]<=26'd1961108; ROM2[9013]<=26'd11120398; ROM3[9013]<=26'd9724858; ROM4[9013]<=26'd23446142;
ROM1[9014]<=26'd1980946; ROM2[9014]<=26'd11129849; ROM3[9014]<=26'd9729126; ROM4[9014]<=26'd23452330;
ROM1[9015]<=26'd1988861; ROM2[9015]<=26'd11132544; ROM3[9015]<=26'd9727300; ROM4[9015]<=26'd23453672;
ROM1[9016]<=26'd1981460; ROM2[9016]<=26'd11130965; ROM3[9016]<=26'd9725041; ROM4[9016]<=26'd23452301;
ROM1[9017]<=26'd1974242; ROM2[9017]<=26'd11132698; ROM3[9017]<=26'd9728537; ROM4[9017]<=26'd23455784;
ROM1[9018]<=26'd1966262; ROM2[9018]<=26'd11130746; ROM3[9018]<=26'd9729231; ROM4[9018]<=26'd23455861;
ROM1[9019]<=26'd1955748; ROM2[9019]<=26'd11125169; ROM3[9019]<=26'd9728202; ROM4[9019]<=26'd23452182;
ROM1[9020]<=26'd1950752; ROM2[9020]<=26'd11120299; ROM3[9020]<=26'd9725980; ROM4[9020]<=26'd23450216;
ROM1[9021]<=26'd1951180; ROM2[9021]<=26'd11118205; ROM3[9021]<=26'd9719774; ROM4[9021]<=26'd23445528;
ROM1[9022]<=26'd1960164; ROM2[9022]<=26'd11115916; ROM3[9022]<=26'd9711319; ROM4[9022]<=26'd23440637;
ROM1[9023]<=26'd1968526; ROM2[9023]<=26'd11114602; ROM3[9023]<=26'd9704404; ROM4[9023]<=26'd23440154;
ROM1[9024]<=26'd1966780; ROM2[9024]<=26'd11116545; ROM3[9024]<=26'd9705567; ROM4[9024]<=26'd23441410;
ROM1[9025]<=26'd1963070; ROM2[9025]<=26'd11118146; ROM3[9025]<=26'd9710605; ROM4[9025]<=26'd23444818;
ROM1[9026]<=26'd1958137; ROM2[9026]<=26'd11117706; ROM3[9026]<=26'd9713657; ROM4[9026]<=26'd23446082;
ROM1[9027]<=26'd1952916; ROM2[9027]<=26'd11117362; ROM3[9027]<=26'd9714451; ROM4[9027]<=26'd23444181;
ROM1[9028]<=26'd1949992; ROM2[9028]<=26'd11118090; ROM3[9028]<=26'd9715478; ROM4[9028]<=26'd23443889;
ROM1[9029]<=26'd1955702; ROM2[9029]<=26'd11121619; ROM3[9029]<=26'd9718336; ROM4[9029]<=26'd23447965;
ROM1[9030]<=26'd1971568; ROM2[9030]<=26'd11129319; ROM3[9030]<=26'd9721324; ROM4[9030]<=26'd23454047;
ROM1[9031]<=26'd1987613; ROM2[9031]<=26'd11135203; ROM3[9031]<=26'd9720199; ROM4[9031]<=26'd23457406;
ROM1[9032]<=26'd1983961; ROM2[9032]<=26'd11129669; ROM3[9032]<=26'd9712711; ROM4[9032]<=26'd23451635;
ROM1[9033]<=26'd1971356; ROM2[9033]<=26'd11121210; ROM3[9033]<=26'd9707440; ROM4[9033]<=26'd23443107;
ROM1[9034]<=26'd1961455; ROM2[9034]<=26'd11116620; ROM3[9034]<=26'd9707905; ROM4[9034]<=26'd23438457;
ROM1[9035]<=26'd1960044; ROM2[9035]<=26'd11119652; ROM3[9035]<=26'd9714903; ROM4[9035]<=26'd23442113;
ROM1[9036]<=26'd1962933; ROM2[9036]<=26'd11128140; ROM3[9036]<=26'd9726759; ROM4[9036]<=26'd23450741;
ROM1[9037]<=26'd1957049; ROM2[9037]<=26'd11123295; ROM3[9037]<=26'd9720749; ROM4[9037]<=26'd23444515;
ROM1[9038]<=26'd1953395; ROM2[9038]<=26'd11115445; ROM3[9038]<=26'd9707804; ROM4[9038]<=26'd23434037;
ROM1[9039]<=26'd1961592; ROM2[9039]<=26'd11112899; ROM3[9039]<=26'd9699304; ROM4[9039]<=26'd23429548;
ROM1[9040]<=26'd1967458; ROM2[9040]<=26'd11112659; ROM3[9040]<=26'd9697396; ROM4[9040]<=26'd23428910;
ROM1[9041]<=26'd1971688; ROM2[9041]<=26'd11120097; ROM3[9041]<=26'd9709928; ROM4[9041]<=26'd23438606;
ROM1[9042]<=26'd1971783; ROM2[9042]<=26'd11126168; ROM3[9042]<=26'd9721038; ROM4[9042]<=26'd23447515;
ROM1[9043]<=26'd1960546; ROM2[9043]<=26'd11118305; ROM3[9043]<=26'd9717912; ROM4[9043]<=26'd23441406;
ROM1[9044]<=26'd1947737; ROM2[9044]<=26'd11108567; ROM3[9044]<=26'd9713387; ROM4[9044]<=26'd23434320;
ROM1[9045]<=26'd1942884; ROM2[9045]<=26'd11108066; ROM3[9045]<=26'd9713625; ROM4[9045]<=26'd23433795;
ROM1[9046]<=26'd1945315; ROM2[9046]<=26'd11107418; ROM3[9046]<=26'd9711323; ROM4[9046]<=26'd23433667;
ROM1[9047]<=26'd1960602; ROM2[9047]<=26'd11113576; ROM3[9047]<=26'd9712667; ROM4[9047]<=26'd23438859;
ROM1[9048]<=26'd1973459; ROM2[9048]<=26'd11118513; ROM3[9048]<=26'd9713372; ROM4[9048]<=26'd23442694;
ROM1[9049]<=26'd1971731; ROM2[9049]<=26'd11117711; ROM3[9049]<=26'd9714303; ROM4[9049]<=26'd23442125;
ROM1[9050]<=26'd1964874; ROM2[9050]<=26'd11118348; ROM3[9050]<=26'd9714456; ROM4[9050]<=26'd23442472;
ROM1[9051]<=26'd1958157; ROM2[9051]<=26'd11117782; ROM3[9051]<=26'd9714745; ROM4[9051]<=26'd23444151;
ROM1[9052]<=26'd1953546; ROM2[9052]<=26'd11117127; ROM3[9052]<=26'd9715844; ROM4[9052]<=26'd23444024;
ROM1[9053]<=26'd1954155; ROM2[9053]<=26'd11122518; ROM3[9053]<=26'd9721116; ROM4[9053]<=26'd23448977;
ROM1[9054]<=26'd1961166; ROM2[9054]<=26'd11129276; ROM3[9054]<=26'd9722818; ROM4[9054]<=26'd23454242;
ROM1[9055]<=26'd1961569; ROM2[9055]<=26'd11121280; ROM3[9055]<=26'd9708347; ROM4[9055]<=26'd23444571;
ROM1[9056]<=26'd1967674; ROM2[9056]<=26'd11118198; ROM3[9056]<=26'd9696802; ROM4[9056]<=26'd23439296;
ROM1[9057]<=26'd1972738; ROM2[9057]<=26'd11124135; ROM3[9057]<=26'd9696764; ROM4[9057]<=26'd23443478;
ROM1[9058]<=26'd1966585; ROM2[9058]<=26'd11122547; ROM3[9058]<=26'd9699435; ROM4[9058]<=26'd23442525;
ROM1[9059]<=26'd1961512; ROM2[9059]<=26'd11124180; ROM3[9059]<=26'd9703594; ROM4[9059]<=26'd23442827;
ROM1[9060]<=26'd1957439; ROM2[9060]<=26'd11124917; ROM3[9060]<=26'd9704999; ROM4[9060]<=26'd23443770;
ROM1[9061]<=26'd1948310; ROM2[9061]<=26'd11120014; ROM3[9061]<=26'd9704550; ROM4[9061]<=26'd23440736;
ROM1[9062]<=26'd1946816; ROM2[9062]<=26'd11118654; ROM3[9062]<=26'd9703860; ROM4[9062]<=26'd23439113;
ROM1[9063]<=26'd1961126; ROM2[9063]<=26'd11126577; ROM3[9063]<=26'd9708868; ROM4[9063]<=26'd23446241;
ROM1[9064]<=26'd1975128; ROM2[9064]<=26'd11130590; ROM3[9064]<=26'd9706535; ROM4[9064]<=26'd23447917;
ROM1[9065]<=26'd1973717; ROM2[9065]<=26'd11124535; ROM3[9065]<=26'd9696750; ROM4[9065]<=26'd23440832;
ROM1[9066]<=26'd1967606; ROM2[9066]<=26'd11122474; ROM3[9066]<=26'd9699052; ROM4[9066]<=26'd23440032;
ROM1[9067]<=26'd1967707; ROM2[9067]<=26'd11128477; ROM3[9067]<=26'd9713027; ROM4[9067]<=26'd23447424;
ROM1[9068]<=26'd1961449; ROM2[9068]<=26'd11127090; ROM3[9068]<=26'd9716879; ROM4[9068]<=26'd23447411;
ROM1[9069]<=26'd1949106; ROM2[9069]<=26'd11116618; ROM3[9069]<=26'd9714002; ROM4[9069]<=26'd23439038;
ROM1[9070]<=26'd1946241; ROM2[9070]<=26'd11114711; ROM3[9070]<=26'd9716016; ROM4[9070]<=26'd23439195;
ROM1[9071]<=26'd1947276; ROM2[9071]<=26'd11114471; ROM3[9071]<=26'd9712105; ROM4[9071]<=26'd23436998;
ROM1[9072]<=26'd1960928; ROM2[9072]<=26'd11116806; ROM3[9072]<=26'd9711594; ROM4[9072]<=26'd23438624;
ROM1[9073]<=26'd1975794; ROM2[9073]<=26'd11123900; ROM3[9073]<=26'd9716005; ROM4[9073]<=26'd23445761;
ROM1[9074]<=26'd1969722; ROM2[9074]<=26'd11119437; ROM3[9074]<=26'd9714030; ROM4[9074]<=26'd23442149;
ROM1[9075]<=26'd1960324; ROM2[9075]<=26'd11112627; ROM3[9075]<=26'd9713227; ROM4[9075]<=26'd23438638;
ROM1[9076]<=26'd1956886; ROM2[9076]<=26'd11111988; ROM3[9076]<=26'd9719879; ROM4[9076]<=26'd23441603;
ROM1[9077]<=26'd1953468; ROM2[9077]<=26'd11113700; ROM3[9077]<=26'd9723921; ROM4[9077]<=26'd23443357;
ROM1[9078]<=26'd1946820; ROM2[9078]<=26'd11113325; ROM3[9078]<=26'd9726917; ROM4[9078]<=26'd23444360;
ROM1[9079]<=26'd1949333; ROM2[9079]<=26'd11113948; ROM3[9079]<=26'd9727907; ROM4[9079]<=26'd23446597;
ROM1[9080]<=26'd1962326; ROM2[9080]<=26'd11117988; ROM3[9080]<=26'd9725732; ROM4[9080]<=26'd23447802;
ROM1[9081]<=26'd1979027; ROM2[9081]<=26'd11121040; ROM3[9081]<=26'd9724200; ROM4[9081]<=26'd23450846;
ROM1[9082]<=26'd1984090; ROM2[9082]<=26'd11123202; ROM3[9082]<=26'd9725340; ROM4[9082]<=26'd23453435;
ROM1[9083]<=26'd1976300; ROM2[9083]<=26'd11122942; ROM3[9083]<=26'd9726199; ROM4[9083]<=26'd23453229;
ROM1[9084]<=26'd1967316; ROM2[9084]<=26'd11122074; ROM3[9084]<=26'd9726856; ROM4[9084]<=26'd23454245;
ROM1[9085]<=26'd1964080; ROM2[9085]<=26'd11123197; ROM3[9085]<=26'd9729366; ROM4[9085]<=26'd23456236;
ROM1[9086]<=26'd1960088; ROM2[9086]<=26'd11124568; ROM3[9086]<=26'd9729696; ROM4[9086]<=26'd23456186;
ROM1[9087]<=26'd1960996; ROM2[9087]<=26'd11125980; ROM3[9087]<=26'd9728351; ROM4[9087]<=26'd23456168;
ROM1[9088]<=26'd1969032; ROM2[9088]<=26'd11128128; ROM3[9088]<=26'd9726103; ROM4[9088]<=26'd23456263;
ROM1[9089]<=26'd1979418; ROM2[9089]<=26'd11129259; ROM3[9089]<=26'd9715416; ROM4[9089]<=26'd23452697;
ROM1[9090]<=26'd1981789; ROM2[9090]<=26'd11126042; ROM3[9090]<=26'd9705816; ROM4[9090]<=26'd23446810;
ROM1[9091]<=26'd1979461; ROM2[9091]<=26'd11126721; ROM3[9091]<=26'd9708934; ROM4[9091]<=26'd23447043;
ROM1[9092]<=26'd1982804; ROM2[9092]<=26'd11139157; ROM3[9092]<=26'd9723141; ROM4[9092]<=26'd23458719;
ROM1[9093]<=26'd1974792; ROM2[9093]<=26'd11139212; ROM3[9093]<=26'd9724435; ROM4[9093]<=26'd23457563;
ROM1[9094]<=26'd1957872; ROM2[9094]<=26'd11127532; ROM3[9094]<=26'd9716388; ROM4[9094]<=26'd23447330;
ROM1[9095]<=26'd1961160; ROM2[9095]<=26'd11133262; ROM3[9095]<=26'd9724526; ROM4[9095]<=26'd23453802;
ROM1[9096]<=26'd1965100; ROM2[9096]<=26'd11133994; ROM3[9096]<=26'd9721191; ROM4[9096]<=26'd23453582;
ROM1[9097]<=26'd1966655; ROM2[9097]<=26'd11124710; ROM3[9097]<=26'd9708479; ROM4[9097]<=26'd23444629;
ROM1[9098]<=26'd1974422; ROM2[9098]<=26'd11125148; ROM3[9098]<=26'd9703070; ROM4[9098]<=26'd23443893;
ROM1[9099]<=26'd1967461; ROM2[9099]<=26'd11120895; ROM3[9099]<=26'd9696249; ROM4[9099]<=26'd23439627;
ROM1[9100]<=26'd1955365; ROM2[9100]<=26'd11113759; ROM3[9100]<=26'd9696186; ROM4[9100]<=26'd23434952;
ROM1[9101]<=26'd1953608; ROM2[9101]<=26'd11116849; ROM3[9101]<=26'd9705484; ROM4[9101]<=26'd23440609;
ROM1[9102]<=26'd1954985; ROM2[9102]<=26'd11122219; ROM3[9102]<=26'd9713882; ROM4[9102]<=26'd23448035;
ROM1[9103]<=26'd1948959; ROM2[9103]<=26'd11121159; ROM3[9103]<=26'd9715642; ROM4[9103]<=26'd23449552;
ROM1[9104]<=26'd1952349; ROM2[9104]<=26'd11124707; ROM3[9104]<=26'd9716756; ROM4[9104]<=26'd23453021;
ROM1[9105]<=26'd1962366; ROM2[9105]<=26'd11125934; ROM3[9105]<=26'd9713100; ROM4[9105]<=26'd23452516;
ROM1[9106]<=26'd1968024; ROM2[9106]<=26'd11118733; ROM3[9106]<=26'd9701821; ROM4[9106]<=26'd23443997;
ROM1[9107]<=26'd1965933; ROM2[9107]<=26'd11115391; ROM3[9107]<=26'd9696071; ROM4[9107]<=26'd23438266;
ROM1[9108]<=26'd1957249; ROM2[9108]<=26'd11113511; ROM3[9108]<=26'd9694342; ROM4[9108]<=26'd23435484;
ROM1[9109]<=26'd1952250; ROM2[9109]<=26'd11114247; ROM3[9109]<=26'd9699271; ROM4[9109]<=26'd23436775;
ROM1[9110]<=26'd1951139; ROM2[9110]<=26'd11116968; ROM3[9110]<=26'd9708351; ROM4[9110]<=26'd23440355;
ROM1[9111]<=26'd1945671; ROM2[9111]<=26'd11114724; ROM3[9111]<=26'd9712131; ROM4[9111]<=26'd23440241;
ROM1[9112]<=26'd1943860; ROM2[9112]<=26'd11110758; ROM3[9112]<=26'd9710734; ROM4[9112]<=26'd23438589;
ROM1[9113]<=26'd1951897; ROM2[9113]<=26'd11111794; ROM3[9113]<=26'd9709983; ROM4[9113]<=26'd23439041;
ROM1[9114]<=26'd1967462; ROM2[9114]<=26'd11117991; ROM3[9114]<=26'd9710267; ROM4[9114]<=26'd23442187;
ROM1[9115]<=26'd1972737; ROM2[9115]<=26'd11118754; ROM3[9115]<=26'd9708111; ROM4[9115]<=26'd23442006;
ROM1[9116]<=26'd1965483; ROM2[9116]<=26'd11114409; ROM3[9116]<=26'd9706864; ROM4[9116]<=26'd23436181;
ROM1[9117]<=26'd1957392; ROM2[9117]<=26'd11113436; ROM3[9117]<=26'd9708116; ROM4[9117]<=26'd23435383;
ROM1[9118]<=26'd1954927; ROM2[9118]<=26'd11114085; ROM3[9118]<=26'd9710471; ROM4[9118]<=26'd23438245;
ROM1[9119]<=26'd1949622; ROM2[9119]<=26'd11114874; ROM3[9119]<=26'd9712690; ROM4[9119]<=26'd23439533;
ROM1[9120]<=26'd1945976; ROM2[9120]<=26'd11114354; ROM3[9120]<=26'd9714497; ROM4[9120]<=26'd23441075;
ROM1[9121]<=26'd1950699; ROM2[9121]<=26'd11115169; ROM3[9121]<=26'd9716182; ROM4[9121]<=26'd23442915;
ROM1[9122]<=26'd1962385; ROM2[9122]<=26'd11115155; ROM3[9122]<=26'd9711646; ROM4[9122]<=26'd23442405;
ROM1[9123]<=26'd1969979; ROM2[9123]<=26'd11112598; ROM3[9123]<=26'd9704018; ROM4[9123]<=26'd23438118;
ROM1[9124]<=26'd1964555; ROM2[9124]<=26'd11111586; ROM3[9124]<=26'd9701766; ROM4[9124]<=26'd23433635;
ROM1[9125]<=26'd1962013; ROM2[9125]<=26'd11116646; ROM3[9125]<=26'd9706378; ROM4[9125]<=26'd23437768;
ROM1[9126]<=26'd1961932; ROM2[9126]<=26'd11124246; ROM3[9126]<=26'd9711932; ROM4[9126]<=26'd23441555;
ROM1[9127]<=26'd1956298; ROM2[9127]<=26'd11122767; ROM3[9127]<=26'd9712958; ROM4[9127]<=26'd23440486;
ROM1[9128]<=26'd1949735; ROM2[9128]<=26'd11119309; ROM3[9128]<=26'd9712715; ROM4[9128]<=26'd23438069;
ROM1[9129]<=26'd1953223; ROM2[9129]<=26'd11121440; ROM3[9129]<=26'd9713794; ROM4[9129]<=26'd23438235;
ROM1[9130]<=26'd1956763; ROM2[9130]<=26'd11117448; ROM3[9130]<=26'd9705803; ROM4[9130]<=26'd23434079;
ROM1[9131]<=26'd1961152; ROM2[9131]<=26'd11110950; ROM3[9131]<=26'd9692679; ROM4[9131]<=26'd23425519;
ROM1[9132]<=26'd1965201; ROM2[9132]<=26'd11112763; ROM3[9132]<=26'd9691527; ROM4[9132]<=26'd23426854;
ROM1[9133]<=26'd1960869; ROM2[9133]<=26'd11113031; ROM3[9133]<=26'd9694579; ROM4[9133]<=26'd23429363;
ROM1[9134]<=26'd1954363; ROM2[9134]<=26'd11113003; ROM3[9134]<=26'd9700395; ROM4[9134]<=26'd23432289;
ROM1[9135]<=26'd1956057; ROM2[9135]<=26'd11120040; ROM3[9135]<=26'd9708533; ROM4[9135]<=26'd23438841;
ROM1[9136]<=26'd1961414; ROM2[9136]<=26'd11129006; ROM3[9136]<=26'd9719547; ROM4[9136]<=26'd23449073;
ROM1[9137]<=26'd1962845; ROM2[9137]<=26'd11130665; ROM3[9137]<=26'd9722065; ROM4[9137]<=26'd23451285;
ROM1[9138]<=26'd1963723; ROM2[9138]<=26'd11126193; ROM3[9138]<=26'd9716067; ROM4[9138]<=26'd23445800;
ROM1[9139]<=26'd1972340; ROM2[9139]<=26'd11123063; ROM3[9139]<=26'd9707965; ROM4[9139]<=26'd23444129;
ROM1[9140]<=26'd1973480; ROM2[9140]<=26'd11117635; ROM3[9140]<=26'd9700029; ROM4[9140]<=26'd23440517;
ROM1[9141]<=26'd1969937; ROM2[9141]<=26'd11117878; ROM3[9141]<=26'd9701029; ROM4[9141]<=26'd23439073;
ROM1[9142]<=26'd1968974; ROM2[9142]<=26'd11122404; ROM3[9142]<=26'd9710272; ROM4[9142]<=26'd23444941;
ROM1[9143]<=26'd1967126; ROM2[9143]<=26'd11124454; ROM3[9143]<=26'd9720199; ROM4[9143]<=26'd23450589;
ROM1[9144]<=26'd1963314; ROM2[9144]<=26'd11124824; ROM3[9144]<=26'd9724618; ROM4[9144]<=26'd23452996;
ROM1[9145]<=26'd1961101; ROM2[9145]<=26'd11125250; ROM3[9145]<=26'd9726188; ROM4[9145]<=26'd23453544;
ROM1[9146]<=26'd1965431; ROM2[9146]<=26'd11125645; ROM3[9146]<=26'd9725066; ROM4[9146]<=26'd23452701;
ROM1[9147]<=26'd1976165; ROM2[9147]<=26'd11128497; ROM3[9147]<=26'd9721899; ROM4[9147]<=26'd23451811;
ROM1[9148]<=26'd1986660; ROM2[9148]<=26'd11132971; ROM3[9148]<=26'd9720825; ROM4[9148]<=26'd23453147;
ROM1[9149]<=26'd1975900; ROM2[9149]<=26'd11123696; ROM3[9149]<=26'd9712205; ROM4[9149]<=26'd23445798;
ROM1[9150]<=26'd1963418; ROM2[9150]<=26'd11117406; ROM3[9150]<=26'd9708834; ROM4[9150]<=26'd23441234;
ROM1[9151]<=26'd1957208; ROM2[9151]<=26'd11116052; ROM3[9151]<=26'd9712030; ROM4[9151]<=26'd23441474;
ROM1[9152]<=26'd1948514; ROM2[9152]<=26'd11112768; ROM3[9152]<=26'd9710336; ROM4[9152]<=26'd23438757;
ROM1[9153]<=26'd1947825; ROM2[9153]<=26'd11115672; ROM3[9153]<=26'd9716729; ROM4[9153]<=26'd23443021;
ROM1[9154]<=26'd1954719; ROM2[9154]<=26'd11119454; ROM3[9154]<=26'd9719377; ROM4[9154]<=26'd23446689;
ROM1[9155]<=26'd1964456; ROM2[9155]<=26'd11120073; ROM3[9155]<=26'd9712697; ROM4[9155]<=26'd23444416;
ROM1[9156]<=26'd1973999; ROM2[9156]<=26'd11118933; ROM3[9156]<=26'd9705525; ROM4[9156]<=26'd23441421;
ROM1[9157]<=26'd1973614; ROM2[9157]<=26'd11118481; ROM3[9157]<=26'd9701882; ROM4[9157]<=26'd23439728;
ROM1[9158]<=26'd1967945; ROM2[9158]<=26'd11118848; ROM3[9158]<=26'd9704368; ROM4[9158]<=26'd23441582;
ROM1[9159]<=26'd1962738; ROM2[9159]<=26'd11117652; ROM3[9159]<=26'd9709324; ROM4[9159]<=26'd23442027;
ROM1[9160]<=26'd1958039; ROM2[9160]<=26'd11115204; ROM3[9160]<=26'd9711897; ROM4[9160]<=26'd23442502;
ROM1[9161]<=26'd1954489; ROM2[9161]<=26'd11116027; ROM3[9161]<=26'd9716464; ROM4[9161]<=26'd23444224;
ROM1[9162]<=26'd1957225; ROM2[9162]<=26'd11119520; ROM3[9162]<=26'd9718696; ROM4[9162]<=26'd23445769;
ROM1[9163]<=26'd1964027; ROM2[9163]<=26'd11120532; ROM3[9163]<=26'd9714849; ROM4[9163]<=26'd23444767;
ROM1[9164]<=26'd1971474; ROM2[9164]<=26'd11118905; ROM3[9164]<=26'd9706593; ROM4[9164]<=26'd23439136;
ROM1[9165]<=26'd1973491; ROM2[9165]<=26'd11115935; ROM3[9165]<=26'd9700464; ROM4[9165]<=26'd23435485;
ROM1[9166]<=26'd1968196; ROM2[9166]<=26'd11114004; ROM3[9166]<=26'd9700912; ROM4[9166]<=26'd23433186;
ROM1[9167]<=26'd1958422; ROM2[9167]<=26'd11112612; ROM3[9167]<=26'd9704417; ROM4[9167]<=26'd23433286;
ROM1[9168]<=26'd1953422; ROM2[9168]<=26'd11112505; ROM3[9168]<=26'd9706345; ROM4[9168]<=26'd23433270;
ROM1[9169]<=26'd1946894; ROM2[9169]<=26'd11111256; ROM3[9169]<=26'd9707417; ROM4[9169]<=26'd23430634;
ROM1[9170]<=26'd1950004; ROM2[9170]<=26'd11119748; ROM3[9170]<=26'd9715904; ROM4[9170]<=26'd23439267;
ROM1[9171]<=26'd1961448; ROM2[9171]<=26'd11127525; ROM3[9171]<=26'd9718549; ROM4[9171]<=26'd23446565;
ROM1[9172]<=26'd1965329; ROM2[9172]<=26'd11121423; ROM3[9172]<=26'd9708800; ROM4[9172]<=26'd23439464;
ROM1[9173]<=26'd1967850; ROM2[9173]<=26'd11117402; ROM3[9173]<=26'd9699051; ROM4[9173]<=26'd23434547;
ROM1[9174]<=26'd1959700; ROM2[9174]<=26'd11109752; ROM3[9174]<=26'd9692905; ROM4[9174]<=26'd23428336;
ROM1[9175]<=26'd1949685; ROM2[9175]<=26'd11105996; ROM3[9175]<=26'd9693345; ROM4[9175]<=26'd23424762;
ROM1[9176]<=26'd1948829; ROM2[9176]<=26'd11109981; ROM3[9176]<=26'd9699264; ROM4[9176]<=26'd23428893;
ROM1[9177]<=26'd1945609; ROM2[9177]<=26'd11109890; ROM3[9177]<=26'd9702856; ROM4[9177]<=26'd23429310;
ROM1[9178]<=26'd1940393; ROM2[9178]<=26'd11108291; ROM3[9178]<=26'd9703898; ROM4[9178]<=26'd23428999;
ROM1[9179]<=26'd1949678; ROM2[9179]<=26'd11114723; ROM3[9179]<=26'd9710226; ROM4[9179]<=26'd23436013;
ROM1[9180]<=26'd1962392; ROM2[9180]<=26'd11116891; ROM3[9180]<=26'd9709061; ROM4[9180]<=26'd23438045;
ROM1[9181]<=26'd1973033; ROM2[9181]<=26'd11115300; ROM3[9181]<=26'd9700909; ROM4[9181]<=26'd23435588;
ROM1[9182]<=26'd1979083; ROM2[9182]<=26'd11119562; ROM3[9182]<=26'd9703958; ROM4[9182]<=26'd23438448;
ROM1[9183]<=26'd1963107; ROM2[9183]<=26'd11109682; ROM3[9183]<=26'd9697699; ROM4[9183]<=26'd23428301;
ROM1[9184]<=26'd1950265; ROM2[9184]<=26'd11103556; ROM3[9184]<=26'd9696103; ROM4[9184]<=26'd23423680;
ROM1[9185]<=26'd1949790; ROM2[9185]<=26'd11107488; ROM3[9185]<=26'd9702818; ROM4[9185]<=26'd23428370;
ROM1[9186]<=26'd1937884; ROM2[9186]<=26'd11101613; ROM3[9186]<=26'd9698551; ROM4[9186]<=26'd23423312;
ROM1[9187]<=26'd1937473; ROM2[9187]<=26'd11102302; ROM3[9187]<=26'd9699294; ROM4[9187]<=26'd23424562;
ROM1[9188]<=26'd1949795; ROM2[9188]<=26'd11109662; ROM3[9188]<=26'd9702556; ROM4[9188]<=26'd23428039;
ROM1[9189]<=26'd1961856; ROM2[9189]<=26'd11111216; ROM3[9189]<=26'd9697001; ROM4[9189]<=26'd23428531;
ROM1[9190]<=26'd1966531; ROM2[9190]<=26'd11111483; ROM3[9190]<=26'd9693311; ROM4[9190]<=26'd23427933;
ROM1[9191]<=26'd1962061; ROM2[9191]<=26'd11110686; ROM3[9191]<=26'd9694502; ROM4[9191]<=26'd23426488;
ROM1[9192]<=26'd1958618; ROM2[9192]<=26'd11113866; ROM3[9192]<=26'd9701803; ROM4[9192]<=26'd23432435;
ROM1[9193]<=26'd1956537; ROM2[9193]<=26'd11118602; ROM3[9193]<=26'd9710091; ROM4[9193]<=26'd23438541;
ROM1[9194]<=26'd1950120; ROM2[9194]<=26'd11116526; ROM3[9194]<=26'd9712347; ROM4[9194]<=26'd23436634;
ROM1[9195]<=26'd1948019; ROM2[9195]<=26'd11115333; ROM3[9195]<=26'd9710979; ROM4[9195]<=26'd23436318;
ROM1[9196]<=26'd1951104; ROM2[9196]<=26'd11114628; ROM3[9196]<=26'd9706298; ROM4[9196]<=26'd23434394;
ROM1[9197]<=26'd1960502; ROM2[9197]<=26'd11114544; ROM3[9197]<=26'd9701147; ROM4[9197]<=26'd23432142;
ROM1[9198]<=26'd1969081; ROM2[9198]<=26'd11114703; ROM3[9198]<=26'd9696579; ROM4[9198]<=26'd23433203;
ROM1[9199]<=26'd1968012; ROM2[9199]<=26'd11115848; ROM3[9199]<=26'd9699136; ROM4[9199]<=26'd23435837;
ROM1[9200]<=26'd1964456; ROM2[9200]<=26'd11118184; ROM3[9200]<=26'd9703848; ROM4[9200]<=26'd23438445;
ROM1[9201]<=26'd1960636; ROM2[9201]<=26'd11118571; ROM3[9201]<=26'd9709118; ROM4[9201]<=26'd23439904;
ROM1[9202]<=26'd1958783; ROM2[9202]<=26'd11121092; ROM3[9202]<=26'd9714422; ROM4[9202]<=26'd23444064;
ROM1[9203]<=26'd1955208; ROM2[9203]<=26'd11121426; ROM3[9203]<=26'd9717083; ROM4[9203]<=26'd23445207;
ROM1[9204]<=26'd1956270; ROM2[9204]<=26'd11119741; ROM3[9204]<=26'd9717529; ROM4[9204]<=26'd23446307;
ROM1[9205]<=26'd1966440; ROM2[9205]<=26'd11122115; ROM3[9205]<=26'd9713613; ROM4[9205]<=26'd23447085;
ROM1[9206]<=26'd1979690; ROM2[9206]<=26'd11124829; ROM3[9206]<=26'd9710549; ROM4[9206]<=26'd23447139;
ROM1[9207]<=26'd1982769; ROM2[9207]<=26'd11126673; ROM3[9207]<=26'd9713169; ROM4[9207]<=26'd23449642;
ROM1[9208]<=26'd1974901; ROM2[9208]<=26'd11126212; ROM3[9208]<=26'd9716716; ROM4[9208]<=26'd23449104;
ROM1[9209]<=26'd1972344; ROM2[9209]<=26'd11129371; ROM3[9209]<=26'd9725551; ROM4[9209]<=26'd23453850;
ROM1[9210]<=26'd1970124; ROM2[9210]<=26'd11132337; ROM3[9210]<=26'd9731719; ROM4[9210]<=26'd23457411;
ROM1[9211]<=26'd1955743; ROM2[9211]<=26'd11121899; ROM3[9211]<=26'd9727427; ROM4[9211]<=26'd23449965;
ROM1[9212]<=26'd1952390; ROM2[9212]<=26'd11118119; ROM3[9212]<=26'd9724630; ROM4[9212]<=26'd23446848;
ROM1[9213]<=26'd1961859; ROM2[9213]<=26'd11121578; ROM3[9213]<=26'd9723180; ROM4[9213]<=26'd23448893;
ROM1[9214]<=26'd1974304; ROM2[9214]<=26'd11122106; ROM3[9214]<=26'd9719399; ROM4[9214]<=26'd23448547;
ROM1[9215]<=26'd1980211; ROM2[9215]<=26'd11124054; ROM3[9215]<=26'd9720315; ROM4[9215]<=26'd23451288;
ROM1[9216]<=26'd1974603; ROM2[9216]<=26'd11121948; ROM3[9216]<=26'd9721251; ROM4[9216]<=26'd23450797;
ROM1[9217]<=26'd1965950; ROM2[9217]<=26'd11119412; ROM3[9217]<=26'd9724735; ROM4[9217]<=26'd23450205;
ROM1[9218]<=26'd1958863; ROM2[9218]<=26'd11116278; ROM3[9218]<=26'd9725590; ROM4[9218]<=26'd23449310;
ROM1[9219]<=26'd1953377; ROM2[9219]<=26'd11113734; ROM3[9219]<=26'd9724459; ROM4[9219]<=26'd23446926;
ROM1[9220]<=26'd1952425; ROM2[9220]<=26'd11114092; ROM3[9220]<=26'd9725732; ROM4[9220]<=26'd23447461;
ROM1[9221]<=26'd1953615; ROM2[9221]<=26'd11112105; ROM3[9221]<=26'd9720531; ROM4[9221]<=26'd23444315;
ROM1[9222]<=26'd1963397; ROM2[9222]<=26'd11111458; ROM3[9222]<=26'd9713938; ROM4[9222]<=26'd23441959;
ROM1[9223]<=26'd1975246; ROM2[9223]<=26'd11116629; ROM3[9223]<=26'd9712589; ROM4[9223]<=26'd23445351;
ROM1[9224]<=26'd1976727; ROM2[9224]<=26'd11120569; ROM3[9224]<=26'd9716213; ROM4[9224]<=26'd23448499;
ROM1[9225]<=26'd1965207; ROM2[9225]<=26'd11113972; ROM3[9225]<=26'd9714210; ROM4[9225]<=26'd23444339;
ROM1[9226]<=26'd1951054; ROM2[9226]<=26'd11107687; ROM3[9226]<=26'd9712112; ROM4[9226]<=26'd23439666;
ROM1[9227]<=26'd1944409; ROM2[9227]<=26'd11107338; ROM3[9227]<=26'd9713694; ROM4[9227]<=26'd23437419;
ROM1[9228]<=26'd1938793; ROM2[9228]<=26'd11105421; ROM3[9228]<=26'd9712398; ROM4[9228]<=26'd23436259;
ROM1[9229]<=26'd1942576; ROM2[9229]<=26'd11110783; ROM3[9229]<=26'd9714278; ROM4[9229]<=26'd23440933;
ROM1[9230]<=26'd1958096; ROM2[9230]<=26'd11119237; ROM3[9230]<=26'd9716935; ROM4[9230]<=26'd23446968;
ROM1[9231]<=26'd1969302; ROM2[9231]<=26'd11118743; ROM3[9231]<=26'd9709257; ROM4[9231]<=26'd23444547;
ROM1[9232]<=26'd1970933; ROM2[9232]<=26'd11119280; ROM3[9232]<=26'd9709444; ROM4[9232]<=26'd23445125;
ROM1[9233]<=26'd1965774; ROM2[9233]<=26'd11118409; ROM3[9233]<=26'd9714033; ROM4[9233]<=26'd23445267;
ROM1[9234]<=26'd1953724; ROM2[9234]<=26'd11113008; ROM3[9234]<=26'd9708619; ROM4[9234]<=26'd23438267;
ROM1[9235]<=26'd1952370; ROM2[9235]<=26'd11117075; ROM3[9235]<=26'd9713446; ROM4[9235]<=26'd23442125;
ROM1[9236]<=26'd1943862; ROM2[9236]<=26'd11114354; ROM3[9236]<=26'd9714626; ROM4[9236]<=26'd23440224;
ROM1[9237]<=26'd1938595; ROM2[9237]<=26'd11108325; ROM3[9237]<=26'd9709271; ROM4[9237]<=26'd23434520;
ROM1[9238]<=26'd1947837; ROM2[9238]<=26'd11108598; ROM3[9238]<=26'd9707860; ROM4[9238]<=26'd23435440;
ROM1[9239]<=26'd1957963; ROM2[9239]<=26'd11110255; ROM3[9239]<=26'd9701334; ROM4[9239]<=26'd23434808;
ROM1[9240]<=26'd1960469; ROM2[9240]<=26'd11109832; ROM3[9240]<=26'd9693877; ROM4[9240]<=26'd23430741;
ROM1[9241]<=26'd1951980; ROM2[9241]<=26'd11105712; ROM3[9241]<=26'd9691116; ROM4[9241]<=26'd23425710;
ROM1[9242]<=26'd1945311; ROM2[9242]<=26'd11105571; ROM3[9242]<=26'd9695420; ROM4[9242]<=26'd23424757;
ROM1[9243]<=26'd1944463; ROM2[9243]<=26'd11107389; ROM3[9243]<=26'd9701444; ROM4[9243]<=26'd23428346;
ROM1[9244]<=26'd1941695; ROM2[9244]<=26'd11110341; ROM3[9244]<=26'd9707930; ROM4[9244]<=26'd23432516;
ROM1[9245]<=26'd1941881; ROM2[9245]<=26'd11112226; ROM3[9245]<=26'd9710853; ROM4[9245]<=26'd23434101;
ROM1[9246]<=26'd1947162; ROM2[9246]<=26'd11112692; ROM3[9246]<=26'd9709555; ROM4[9246]<=26'd23435806;
ROM1[9247]<=26'd1959635; ROM2[9247]<=26'd11114280; ROM3[9247]<=26'd9706448; ROM4[9247]<=26'd23435464;
ROM1[9248]<=26'd1974496; ROM2[9248]<=26'd11117964; ROM3[9248]<=26'd9707107; ROM4[9248]<=26'd23440006;
ROM1[9249]<=26'd1968354; ROM2[9249]<=26'd11113561; ROM3[9249]<=26'd9705890; ROM4[9249]<=26'd23437690;
ROM1[9250]<=26'd1956841; ROM2[9250]<=26'd11107203; ROM3[9250]<=26'd9704808; ROM4[9250]<=26'd23433830;
ROM1[9251]<=26'd1950296; ROM2[9251]<=26'd11105468; ROM3[9251]<=26'd9709132; ROM4[9251]<=26'd23434532;
ROM1[9252]<=26'd1944497; ROM2[9252]<=26'd11103513; ROM3[9252]<=26'd9710463; ROM4[9252]<=26'd23432917;
ROM1[9253]<=26'd1944998; ROM2[9253]<=26'd11105472; ROM3[9253]<=26'd9717274; ROM4[9253]<=26'd23438115;
ROM1[9254]<=26'd1950177; ROM2[9254]<=26'd11110378; ROM3[9254]<=26'd9721949; ROM4[9254]<=26'd23442474;
ROM1[9255]<=26'd1956238; ROM2[9255]<=26'd11109541; ROM3[9255]<=26'd9716031; ROM4[9255]<=26'd23439553;
ROM1[9256]<=26'd1965146; ROM2[9256]<=26'd11108441; ROM3[9256]<=26'd9709464; ROM4[9256]<=26'd23436513;
ROM1[9257]<=26'd1967992; ROM2[9257]<=26'd11111612; ROM3[9257]<=26'd9708943; ROM4[9257]<=26'd23438551;
ROM1[9258]<=26'd1967243; ROM2[9258]<=26'd11115258; ROM3[9258]<=26'd9713682; ROM4[9258]<=26'd23442452;
ROM1[9259]<=26'd1965943; ROM2[9259]<=26'd11117511; ROM3[9259]<=26'd9719275; ROM4[9259]<=26'd23445719;
ROM1[9260]<=26'd1959854; ROM2[9260]<=26'd11116260; ROM3[9260]<=26'd9720347; ROM4[9260]<=26'd23447255;
ROM1[9261]<=26'd1950566; ROM2[9261]<=26'd11112573; ROM3[9261]<=26'd9717782; ROM4[9261]<=26'd23441965;
ROM1[9262]<=26'd1951650; ROM2[9262]<=26'd11115158; ROM3[9262]<=26'd9717107; ROM4[9262]<=26'd23443577;
ROM1[9263]<=26'd1960501; ROM2[9263]<=26'd11118926; ROM3[9263]<=26'd9715758; ROM4[9263]<=26'd23447880;
ROM1[9264]<=26'd1976041; ROM2[9264]<=26'd11122159; ROM3[9264]<=26'd9711919; ROM4[9264]<=26'd23449489;
ROM1[9265]<=26'd1985743; ROM2[9265]<=26'd11127563; ROM3[9265]<=26'd9714123; ROM4[9265]<=26'd23455904;
ROM1[9266]<=26'd1973738; ROM2[9266]<=26'd11120918; ROM3[9266]<=26'd9711185; ROM4[9266]<=26'd23451334;
ROM1[9267]<=26'd1960982; ROM2[9267]<=26'd11115337; ROM3[9267]<=26'd9709034; ROM4[9267]<=26'd23446254;
ROM1[9268]<=26'd1957912; ROM2[9268]<=26'd11119297; ROM3[9268]<=26'd9715882; ROM4[9268]<=26'd23450250;
ROM1[9269]<=26'd1954689; ROM2[9269]<=26'd11120077; ROM3[9269]<=26'd9720268; ROM4[9269]<=26'd23451557;
ROM1[9270]<=26'd1951733; ROM2[9270]<=26'd11117853; ROM3[9270]<=26'd9719943; ROM4[9270]<=26'd23449667;
ROM1[9271]<=26'd1952625; ROM2[9271]<=26'd11114322; ROM3[9271]<=26'd9715520; ROM4[9271]<=26'd23445996;
ROM1[9272]<=26'd1959497; ROM2[9272]<=26'd11111029; ROM3[9272]<=26'd9708590; ROM4[9272]<=26'd23440119;
ROM1[9273]<=26'd1967501; ROM2[9273]<=26'd11111541; ROM3[9273]<=26'd9703142; ROM4[9273]<=26'd23438155;
ROM1[9274]<=26'd1970353; ROM2[9274]<=26'd11115907; ROM3[9274]<=26'd9708250; ROM4[9274]<=26'd23441448;
ROM1[9275]<=26'd1967679; ROM2[9275]<=26'd11120511; ROM3[9275]<=26'd9716779; ROM4[9275]<=26'd23444643;
ROM1[9276]<=26'd1960826; ROM2[9276]<=26'd11118462; ROM3[9276]<=26'd9719671; ROM4[9276]<=26'd23445229;
ROM1[9277]<=26'd1951445; ROM2[9277]<=26'd11112422; ROM3[9277]<=26'd9718232; ROM4[9277]<=26'd23442144;
ROM1[9278]<=26'd1944843; ROM2[9278]<=26'd11111562; ROM3[9278]<=26'd9719244; ROM4[9278]<=26'd23440913;
ROM1[9279]<=26'd1944968; ROM2[9279]<=26'd11110083; ROM3[9279]<=26'd9715773; ROM4[9279]<=26'd23438252;
ROM1[9280]<=26'd1950798; ROM2[9280]<=26'd11106583; ROM3[9280]<=26'd9708898; ROM4[9280]<=26'd23434038;
ROM1[9281]<=26'd1961053; ROM2[9281]<=26'd11106094; ROM3[9281]<=26'd9703517; ROM4[9281]<=26'd23432747;
ROM1[9282]<=26'd1960506; ROM2[9282]<=26'd11104146; ROM3[9282]<=26'd9700620; ROM4[9282]<=26'd23430507;
ROM1[9283]<=26'd1956520; ROM2[9283]<=26'd11104471; ROM3[9283]<=26'd9705028; ROM4[9283]<=26'd23432754;
ROM1[9284]<=26'd1949232; ROM2[9284]<=26'd11104960; ROM3[9284]<=26'd9709770; ROM4[9284]<=26'd23434401;
ROM1[9285]<=26'd1945115; ROM2[9285]<=26'd11107028; ROM3[9285]<=26'd9715239; ROM4[9285]<=26'd23435880;
ROM1[9286]<=26'd1940194; ROM2[9286]<=26'd11107521; ROM3[9286]<=26'd9719182; ROM4[9286]<=26'd23439536;
ROM1[9287]<=26'd1937579; ROM2[9287]<=26'd11107344; ROM3[9287]<=26'd9719408; ROM4[9287]<=26'd23440042;
ROM1[9288]<=26'd1950077; ROM2[9288]<=26'd11112433; ROM3[9288]<=26'd9719085; ROM4[9288]<=26'd23442756;
ROM1[9289]<=26'd1965069; ROM2[9289]<=26'd11115053; ROM3[9289]<=26'd9712152; ROM4[9289]<=26'd23442338;
ROM1[9290]<=26'd1971887; ROM2[9290]<=26'd11115305; ROM3[9290]<=26'd9709360; ROM4[9290]<=26'd23440033;
ROM1[9291]<=26'd1973745; ROM2[9291]<=26'd11119594; ROM3[9291]<=26'd9714696; ROM4[9291]<=26'd23444111;
ROM1[9292]<=26'd1968645; ROM2[9292]<=26'd11121056; ROM3[9292]<=26'd9717246; ROM4[9292]<=26'd23445667;
ROM1[9293]<=26'd1960900; ROM2[9293]<=26'd11119284; ROM3[9293]<=26'd9717581; ROM4[9293]<=26'd23444174;
ROM1[9294]<=26'd1948858; ROM2[9294]<=26'd11113096; ROM3[9294]<=26'd9712026; ROM4[9294]<=26'd23436955;
ROM1[9295]<=26'd1937969; ROM2[9295]<=26'd11104154; ROM3[9295]<=26'd9702543; ROM4[9295]<=26'd23426182;
ROM1[9296]<=26'd1940690; ROM2[9296]<=26'd11102199; ROM3[9296]<=26'd9696485; ROM4[9296]<=26'd23421061;
ROM1[9297]<=26'd1956607; ROM2[9297]<=26'd11106918; ROM3[9297]<=26'd9694038; ROM4[9297]<=26'd23423197;
ROM1[9298]<=26'd1967876; ROM2[9298]<=26'd11110096; ROM3[9298]<=26'd9692662; ROM4[9298]<=26'd23426040;
ROM1[9299]<=26'd1969195; ROM2[9299]<=26'd11115004; ROM3[9299]<=26'd9696417; ROM4[9299]<=26'd23430747;
ROM1[9300]<=26'd1968439; ROM2[9300]<=26'd11122020; ROM3[9300]<=26'd9704568; ROM4[9300]<=26'd23438317;
ROM1[9301]<=26'd1955268; ROM2[9301]<=26'd11114811; ROM3[9301]<=26'd9701168; ROM4[9301]<=26'd23432827;
ROM1[9302]<=26'd1948979; ROM2[9302]<=26'd11113492; ROM3[9302]<=26'd9701681; ROM4[9302]<=26'd23431944;
ROM1[9303]<=26'd1949451; ROM2[9303]<=26'd11115498; ROM3[9303]<=26'd9709183; ROM4[9303]<=26'd23436236;
ROM1[9304]<=26'd1945821; ROM2[9304]<=26'd11109834; ROM3[9304]<=26'd9703537; ROM4[9304]<=26'd23430829;
ROM1[9305]<=26'd1955180; ROM2[9305]<=26'd11111054; ROM3[9305]<=26'd9699687; ROM4[9305]<=26'd23430554;
ROM1[9306]<=26'd1972715; ROM2[9306]<=26'd11117871; ROM3[9306]<=26'd9701470; ROM4[9306]<=26'd23436684;
ROM1[9307]<=26'd1981074; ROM2[9307]<=26'd11126374; ROM3[9307]<=26'd9706352; ROM4[9307]<=26'd23443882;
ROM1[9308]<=26'd1971363; ROM2[9308]<=26'd11121300; ROM3[9308]<=26'd9706448; ROM4[9308]<=26'd23440699;
ROM1[9309]<=26'd1958661; ROM2[9309]<=26'd11114644; ROM3[9309]<=26'd9703994; ROM4[9309]<=26'd23435883;
ROM1[9310]<=26'd1958501; ROM2[9310]<=26'd11118618; ROM3[9310]<=26'd9709990; ROM4[9310]<=26'd23440192;
ROM1[9311]<=26'd1949432; ROM2[9311]<=26'd11114170; ROM3[9311]<=26'd9709840; ROM4[9311]<=26'd23436117;
ROM1[9312]<=26'd1946154; ROM2[9312]<=26'd11112426; ROM3[9312]<=26'd9706763; ROM4[9312]<=26'd23433584;
ROM1[9313]<=26'd1959849; ROM2[9313]<=26'd11122000; ROM3[9313]<=26'd9711066; ROM4[9313]<=26'd23439246;
ROM1[9314]<=26'd1970131; ROM2[9314]<=26'd11121558; ROM3[9314]<=26'd9706274; ROM4[9314]<=26'd23436677;
ROM1[9315]<=26'd1967705; ROM2[9315]<=26'd11115853; ROM3[9315]<=26'd9695919; ROM4[9315]<=26'd23430450;
ROM1[9316]<=26'd1962409; ROM2[9316]<=26'd11114679; ROM3[9316]<=26'd9697482; ROM4[9316]<=26'd23430064;
ROM1[9317]<=26'd1957654; ROM2[9317]<=26'd11115577; ROM3[9317]<=26'd9705805; ROM4[9317]<=26'd23433077;
ROM1[9318]<=26'd1951952; ROM2[9318]<=26'd11114716; ROM3[9318]<=26'd9706280; ROM4[9318]<=26'd23432825;
ROM1[9319]<=26'd1944988; ROM2[9319]<=26'd11110670; ROM3[9319]<=26'd9706596; ROM4[9319]<=26'd23430586;
ROM1[9320]<=26'd1943202; ROM2[9320]<=26'd11111995; ROM3[9320]<=26'd9710989; ROM4[9320]<=26'd23433939;
ROM1[9321]<=26'd1949772; ROM2[9321]<=26'd11113509; ROM3[9321]<=26'd9711917; ROM4[9321]<=26'd23437142;
ROM1[9322]<=26'd1963729; ROM2[9322]<=26'd11116470; ROM3[9322]<=26'd9712137; ROM4[9322]<=26'd23439570;
ROM1[9323]<=26'd1967444; ROM2[9323]<=26'd11113077; ROM3[9323]<=26'd9705083; ROM4[9323]<=26'd23436234;
ROM1[9324]<=26'd1961097; ROM2[9324]<=26'd11108420; ROM3[9324]<=26'd9701246; ROM4[9324]<=26'd23432093;
ROM1[9325]<=26'd1955115; ROM2[9325]<=26'd11109690; ROM3[9325]<=26'd9705737; ROM4[9325]<=26'd23434121;
ROM1[9326]<=26'd1946977; ROM2[9326]<=26'd11107857; ROM3[9326]<=26'd9706920; ROM4[9326]<=26'd23432335;
ROM1[9327]<=26'd1942333; ROM2[9327]<=26'd11107811; ROM3[9327]<=26'd9709548; ROM4[9327]<=26'd23432397;
ROM1[9328]<=26'd1940932; ROM2[9328]<=26'd11110358; ROM3[9328]<=26'd9713226; ROM4[9328]<=26'd23436299;
ROM1[9329]<=26'd1944457; ROM2[9329]<=26'd11111846; ROM3[9329]<=26'd9712667; ROM4[9329]<=26'd23436879;
ROM1[9330]<=26'd1954128; ROM2[9330]<=26'd11113617; ROM3[9330]<=26'd9708439; ROM4[9330]<=26'd23436429;
ROM1[9331]<=26'd1967696; ROM2[9331]<=26'd11116641; ROM3[9331]<=26'd9705838; ROM4[9331]<=26'd23438195;
ROM1[9332]<=26'd1973883; ROM2[9332]<=26'd11120930; ROM3[9332]<=26'd9710593; ROM4[9332]<=26'd23442078;
ROM1[9333]<=26'd1969893; ROM2[9333]<=26'd11122579; ROM3[9333]<=26'd9715320; ROM4[9333]<=26'd23444455;
ROM1[9334]<=26'd1956502; ROM2[9334]<=26'd11113776; ROM3[9334]<=26'd9712018; ROM4[9334]<=26'd23438242;
ROM1[9335]<=26'd1953221; ROM2[9335]<=26'd11114331; ROM3[9335]<=26'd9715334; ROM4[9335]<=26'd23440889;
ROM1[9336]<=26'd1948974; ROM2[9336]<=26'd11115484; ROM3[9336]<=26'd9719425; ROM4[9336]<=26'd23443536;
ROM1[9337]<=26'd1947932; ROM2[9337]<=26'd11114117; ROM3[9337]<=26'd9717808; ROM4[9337]<=26'd23442262;
ROM1[9338]<=26'd1963533; ROM2[9338]<=26'd11123636; ROM3[9338]<=26'd9723819; ROM4[9338]<=26'd23450245;
ROM1[9339]<=26'd1981477; ROM2[9339]<=26'd11133007; ROM3[9339]<=26'd9726267; ROM4[9339]<=26'd23455860;
ROM1[9340]<=26'd1981035; ROM2[9340]<=26'd11127493; ROM3[9340]<=26'd9716842; ROM4[9340]<=26'd23449652;
ROM1[9341]<=26'd1967500; ROM2[9341]<=26'd11117587; ROM3[9341]<=26'd9708963; ROM4[9341]<=26'd23439009;
ROM1[9342]<=26'd1959540; ROM2[9342]<=26'd11116814; ROM3[9342]<=26'd9711734; ROM4[9342]<=26'd23437641;
ROM1[9343]<=26'd1957596; ROM2[9343]<=26'd11119002; ROM3[9343]<=26'd9717332; ROM4[9343]<=26'd23442321;
ROM1[9344]<=26'd1958951; ROM2[9344]<=26'd11125490; ROM3[9344]<=26'd9725968; ROM4[9344]<=26'd23447597;
ROM1[9345]<=26'd1954430; ROM2[9345]<=26'd11122604; ROM3[9345]<=26'd9725000; ROM4[9345]<=26'd23445715;
ROM1[9346]<=26'd1952584; ROM2[9346]<=26'd11114448; ROM3[9346]<=26'd9717184; ROM4[9346]<=26'd23439857;
ROM1[9347]<=26'd1960714; ROM2[9347]<=26'd11112881; ROM3[9347]<=26'd9709626; ROM4[9347]<=26'd23434949;
ROM1[9348]<=26'd1972309; ROM2[9348]<=26'd11117644; ROM3[9348]<=26'd9707643; ROM4[9348]<=26'd23438356;
ROM1[9349]<=26'd1976816; ROM2[9349]<=26'd11125063; ROM3[9349]<=26'd9714749; ROM4[9349]<=26'd23446194;
ROM1[9350]<=26'd1974534; ROM2[9350]<=26'd11129004; ROM3[9350]<=26'd9721247; ROM4[9350]<=26'd23450906;
ROM1[9351]<=26'd1967435; ROM2[9351]<=26'd11127414; ROM3[9351]<=26'd9724717; ROM4[9351]<=26'd23451344;
ROM1[9352]<=26'd1960331; ROM2[9352]<=26'd11124264; ROM3[9352]<=26'd9726171; ROM4[9352]<=26'd23450246;
ROM1[9353]<=26'd1951485; ROM2[9353]<=26'd11118971; ROM3[9353]<=26'd9723239; ROM4[9353]<=26'd23446850;
ROM1[9354]<=26'd1950138; ROM2[9354]<=26'd11117936; ROM3[9354]<=26'd9718538; ROM4[9354]<=26'd23443273;
ROM1[9355]<=26'd1957909; ROM2[9355]<=26'd11116945; ROM3[9355]<=26'd9712176; ROM4[9355]<=26'd23440290;
ROM1[9356]<=26'd1968087; ROM2[9356]<=26'd11116502; ROM3[9356]<=26'd9705462; ROM4[9356]<=26'd23437156;
ROM1[9357]<=26'd1977028; ROM2[9357]<=26'd11123210; ROM3[9357]<=26'd9712377; ROM4[9357]<=26'd23444840;
ROM1[9358]<=26'd1971457; ROM2[9358]<=26'd11126110; ROM3[9358]<=26'd9716928; ROM4[9358]<=26'd23448989;
ROM1[9359]<=26'd1960724; ROM2[9359]<=26'd11125173; ROM3[9359]<=26'd9717489; ROM4[9359]<=26'd23446864;
ROM1[9360]<=26'd1954027; ROM2[9360]<=26'd11123101; ROM3[9360]<=26'd9719031; ROM4[9360]<=26'd23447319;
ROM1[9361]<=26'd1945320; ROM2[9361]<=26'd11119798; ROM3[9361]<=26'd9717130; ROM4[9361]<=26'd23442365;
ROM1[9362]<=26'd1947787; ROM2[9362]<=26'd11121852; ROM3[9362]<=26'd9718284; ROM4[9362]<=26'd23443254;
ROM1[9363]<=26'd1959642; ROM2[9363]<=26'd11125130; ROM3[9363]<=26'd9717390; ROM4[9363]<=26'd23446440;
ROM1[9364]<=26'd1972167; ROM2[9364]<=26'd11124883; ROM3[9364]<=26'd9710834; ROM4[9364]<=26'd23442888;
ROM1[9365]<=26'd1976125; ROM2[9365]<=26'd11123202; ROM3[9365]<=26'd9705611; ROM4[9365]<=26'd23441529;
ROM1[9366]<=26'd1969300; ROM2[9366]<=26'd11120350; ROM3[9366]<=26'd9703527; ROM4[9366]<=26'd23437738;
ROM1[9367]<=26'd1960494; ROM2[9367]<=26'd11117586; ROM3[9367]<=26'd9703661; ROM4[9367]<=26'd23434043;
ROM1[9368]<=26'd1956940; ROM2[9368]<=26'd11117962; ROM3[9368]<=26'd9706348; ROM4[9368]<=26'd23435501;
ROM1[9369]<=26'd1952608; ROM2[9369]<=26'd11118656; ROM3[9369]<=26'd9710387; ROM4[9369]<=26'd23435706;
ROM1[9370]<=26'd1950769; ROM2[9370]<=26'd11119580; ROM3[9370]<=26'd9711782; ROM4[9370]<=26'd23436115;
ROM1[9371]<=26'd1951970; ROM2[9371]<=26'd11116169; ROM3[9371]<=26'd9706104; ROM4[9371]<=26'd23433344;
ROM1[9372]<=26'd1957898; ROM2[9372]<=26'd11111965; ROM3[9372]<=26'd9695327; ROM4[9372]<=26'd23427107;
ROM1[9373]<=26'd1962242; ROM2[9373]<=26'd11111174; ROM3[9373]<=26'd9687030; ROM4[9373]<=26'd23424206;
ROM1[9374]<=26'd1958080; ROM2[9374]<=26'd11109827; ROM3[9374]<=26'd9686885; ROM4[9374]<=26'd23423950;
ROM1[9375]<=26'd1954604; ROM2[9375]<=26'd11112511; ROM3[9375]<=26'd9692436; ROM4[9375]<=26'd23426984;
ROM1[9376]<=26'd1947596; ROM2[9376]<=26'd11110406; ROM3[9376]<=26'd9695348; ROM4[9376]<=26'd23427888;
ROM1[9377]<=26'd1944029; ROM2[9377]<=26'd11110356; ROM3[9377]<=26'd9702172; ROM4[9377]<=26'd23431528;
ROM1[9378]<=26'd1938811; ROM2[9378]<=26'd11108076; ROM3[9378]<=26'd9705218; ROM4[9378]<=26'd23431421;
ROM1[9379]<=26'd1938528; ROM2[9379]<=26'd11105493; ROM3[9379]<=26'd9704916; ROM4[9379]<=26'd23429444;
ROM1[9380]<=26'd1951375; ROM2[9380]<=26'd11111758; ROM3[9380]<=26'd9706298; ROM4[9380]<=26'd23433160;
ROM1[9381]<=26'd1960666; ROM2[9381]<=26'd11111650; ROM3[9381]<=26'd9699088; ROM4[9381]<=26'd23431032;
ROM1[9382]<=26'd1949759; ROM2[9382]<=26'd11099560; ROM3[9382]<=26'd9687523; ROM4[9382]<=26'd23419912;
ROM1[9383]<=26'd1938648; ROM2[9383]<=26'd11093634; ROM3[9383]<=26'd9687860; ROM4[9383]<=26'd23415445;
ROM1[9384]<=26'd1938865; ROM2[9384]<=26'd11100828; ROM3[9384]<=26'd9702323; ROM4[9384]<=26'd23422818;
ROM1[9385]<=26'd1941354; ROM2[9385]<=26'd11108394; ROM3[9385]<=26'd9713318; ROM4[9385]<=26'd23430176;
ROM1[9386]<=26'd1946589; ROM2[9386]<=26'd11117688; ROM3[9386]<=26'd9724789; ROM4[9386]<=26'd23440627;
ROM1[9387]<=26'd1954896; ROM2[9387]<=26'd11125043; ROM3[9387]<=26'd9731141; ROM4[9387]<=26'd23447803;
ROM1[9388]<=26'd1960696; ROM2[9388]<=26'd11125114; ROM3[9388]<=26'd9726636; ROM4[9388]<=26'd23445044;
ROM1[9389]<=26'd1972666; ROM2[9389]<=26'd11123987; ROM3[9389]<=26'd9721402; ROM4[9389]<=26'd23443926;
ROM1[9390]<=26'd1976971; ROM2[9390]<=26'd11123295; ROM3[9390]<=26'd9718388; ROM4[9390]<=26'd23442185;
ROM1[9391]<=26'd1971099; ROM2[9391]<=26'd11124027; ROM3[9391]<=26'd9719554; ROM4[9391]<=26'd23442072;
ROM1[9392]<=26'd1970123; ROM2[9392]<=26'd11127644; ROM3[9392]<=26'd9727147; ROM4[9392]<=26'd23449584;
ROM1[9393]<=26'd1965485; ROM2[9393]<=26'd11127024; ROM3[9393]<=26'd9727911; ROM4[9393]<=26'd23448103;
ROM1[9394]<=26'd1958579; ROM2[9394]<=26'd11124114; ROM3[9394]<=26'd9726517; ROM4[9394]<=26'd23445552;
ROM1[9395]<=26'd1957525; ROM2[9395]<=26'd11124333; ROM3[9395]<=26'd9727613; ROM4[9395]<=26'd23447178;
ROM1[9396]<=26'd1964940; ROM2[9396]<=26'd11127826; ROM3[9396]<=26'd9727167; ROM4[9396]<=26'd23451709;
ROM1[9397]<=26'd1972540; ROM2[9397]<=26'd11124143; ROM3[9397]<=26'd9717513; ROM4[9397]<=26'd23448480;
ROM1[9398]<=26'd1978727; ROM2[9398]<=26'd11123373; ROM3[9398]<=26'd9708991; ROM4[9398]<=26'd23444351;
ROM1[9399]<=26'd1976320; ROM2[9399]<=26'd11124061; ROM3[9399]<=26'd9708211; ROM4[9399]<=26'd23444087;
ROM1[9400]<=26'd1961387; ROM2[9400]<=26'd11115110; ROM3[9400]<=26'd9704090; ROM4[9400]<=26'd23434767;
ROM1[9401]<=26'd1953939; ROM2[9401]<=26'd11113682; ROM3[9401]<=26'd9707589; ROM4[9401]<=26'd23432981;
ROM1[9402]<=26'd1950393; ROM2[9402]<=26'd11114317; ROM3[9402]<=26'd9714015; ROM4[9402]<=26'd23436703;
ROM1[9403]<=26'd1943199; ROM2[9403]<=26'd11110284; ROM3[9403]<=26'd9712540; ROM4[9403]<=26'd23433879;
ROM1[9404]<=26'd1946485; ROM2[9404]<=26'd11112858; ROM3[9404]<=26'd9713213; ROM4[9404]<=26'd23433718;
ROM1[9405]<=26'd1957236; ROM2[9405]<=26'd11116970; ROM3[9405]<=26'd9711586; ROM4[9405]<=26'd23435556;
ROM1[9406]<=26'd1967444; ROM2[9406]<=26'd11117936; ROM3[9406]<=26'd9705626; ROM4[9406]<=26'd23434866;
ROM1[9407]<=26'd1969236; ROM2[9407]<=26'd11120480; ROM3[9407]<=26'd9707845; ROM4[9407]<=26'd23437602;
ROM1[9408]<=26'd1966682; ROM2[9408]<=26'd11123633; ROM3[9408]<=26'd9714024; ROM4[9408]<=26'd23441427;
ROM1[9409]<=26'd1960459; ROM2[9409]<=26'd11123539; ROM3[9409]<=26'd9717908; ROM4[9409]<=26'd23442376;
ROM1[9410]<=26'd1954160; ROM2[9410]<=26'd11121648; ROM3[9410]<=26'd9719618; ROM4[9410]<=26'd23443293;
ROM1[9411]<=26'd1948759; ROM2[9411]<=26'd11121082; ROM3[9411]<=26'd9723018; ROM4[9411]<=26'd23443572;
ROM1[9412]<=26'd1944856; ROM2[9412]<=26'd11116587; ROM3[9412]<=26'd9719035; ROM4[9412]<=26'd23438821;
ROM1[9413]<=26'd1953624; ROM2[9413]<=26'd11117819; ROM3[9413]<=26'd9716556; ROM4[9413]<=26'd23439320;
ROM1[9414]<=26'd1971515; ROM2[9414]<=26'd11122234; ROM3[9414]<=26'd9715419; ROM4[9414]<=26'd23441786;
ROM1[9415]<=26'd1981074; ROM2[9415]<=26'd11123266; ROM3[9415]<=26'd9714639; ROM4[9415]<=26'd23443723;
ROM1[9416]<=26'd1980825; ROM2[9416]<=26'd11126122; ROM3[9416]<=26'd9720928; ROM4[9416]<=26'd23448152;
ROM1[9417]<=26'd1972524; ROM2[9417]<=26'd11124045; ROM3[9417]<=26'd9725261; ROM4[9417]<=26'd23447975;
ROM1[9418]<=26'd1966138; ROM2[9418]<=26'd11121531; ROM3[9418]<=26'd9729212; ROM4[9418]<=26'd23447708;
ROM1[9419]<=26'd1962604; ROM2[9419]<=26'd11122851; ROM3[9419]<=26'd9733120; ROM4[9419]<=26'd23449231;
ROM1[9420]<=26'd1955858; ROM2[9420]<=26'd11121150; ROM3[9420]<=26'd9729732; ROM4[9420]<=26'd23446808;
ROM1[9421]<=26'd1957536; ROM2[9421]<=26'd11119203; ROM3[9421]<=26'd9723828; ROM4[9421]<=26'd23443765;
ROM1[9422]<=26'd1967605; ROM2[9422]<=26'd11117909; ROM3[9422]<=26'd9717475; ROM4[9422]<=26'd23440006;
ROM1[9423]<=26'd1969420; ROM2[9423]<=26'd11112794; ROM3[9423]<=26'd9708691; ROM4[9423]<=26'd23434341;
ROM1[9424]<=26'd1961021; ROM2[9424]<=26'd11105634; ROM3[9424]<=26'd9704950; ROM4[9424]<=26'd23428810;
ROM1[9425]<=26'd1955691; ROM2[9425]<=26'd11102986; ROM3[9425]<=26'd9705387; ROM4[9425]<=26'd23427048;
ROM1[9426]<=26'd1956038; ROM2[9426]<=26'd11107308; ROM3[9426]<=26'd9710105; ROM4[9426]<=26'd23430814;
ROM1[9427]<=26'd1950692; ROM2[9427]<=26'd11107805; ROM3[9427]<=26'd9711196; ROM4[9427]<=26'd23429013;
ROM1[9428]<=26'd1941729; ROM2[9428]<=26'd11104708; ROM3[9428]<=26'd9707499; ROM4[9428]<=26'd23424656;
ROM1[9429]<=26'd1944948; ROM2[9429]<=26'd11109715; ROM3[9429]<=26'd9711399; ROM4[9429]<=26'd23427835;
ROM1[9430]<=26'd1955077; ROM2[9430]<=26'd11114426; ROM3[9430]<=26'd9711632; ROM4[9430]<=26'd23429293;
ROM1[9431]<=26'd1962907; ROM2[9431]<=26'd11110280; ROM3[9431]<=26'd9701018; ROM4[9431]<=26'd23424482;
ROM1[9432]<=26'd1968803; ROM2[9432]<=26'd11114007; ROM3[9432]<=26'd9703372; ROM4[9432]<=26'd23428997;
ROM1[9433]<=26'd1971468; ROM2[9433]<=26'd11121105; ROM3[9433]<=26'd9711504; ROM4[9433]<=26'd23437011;
ROM1[9434]<=26'd1968209; ROM2[9434]<=26'd11124833; ROM3[9434]<=26'd9718732; ROM4[9434]<=26'd23442130;
ROM1[9435]<=26'd1970692; ROM2[9435]<=26'd11132885; ROM3[9435]<=26'd9731620; ROM4[9435]<=26'd23452358;
ROM1[9436]<=26'd1957526; ROM2[9436]<=26'd11123349; ROM3[9436]<=26'd9725594; ROM4[9436]<=26'd23442815;
ROM1[9437]<=26'd1942035; ROM2[9437]<=26'd11110801; ROM3[9437]<=26'd9714054; ROM4[9437]<=26'd23428606;
ROM1[9438]<=26'd1944893; ROM2[9438]<=26'd11106129; ROM3[9438]<=26'd9707386; ROM4[9438]<=26'd23425348;
ROM1[9439]<=26'd1956453; ROM2[9439]<=26'd11104898; ROM3[9439]<=26'd9699417; ROM4[9439]<=26'd23423993;
ROM1[9440]<=26'd1963762; ROM2[9440]<=26'd11107094; ROM3[9440]<=26'd9699548; ROM4[9440]<=26'd23425971;
ROM1[9441]<=26'd1961152; ROM2[9441]<=26'd11107272; ROM3[9441]<=26'd9704749; ROM4[9441]<=26'd23429315;
ROM1[9442]<=26'd1954075; ROM2[9442]<=26'd11108359; ROM3[9442]<=26'd9710197; ROM4[9442]<=26'd23432691;
ROM1[9443]<=26'd1950880; ROM2[9443]<=26'd11111087; ROM3[9443]<=26'd9716071; ROM4[9443]<=26'd23435462;
ROM1[9444]<=26'd1953977; ROM2[9444]<=26'd11120125; ROM3[9444]<=26'd9727798; ROM4[9444]<=26'd23445083;
ROM1[9445]<=26'd1950687; ROM2[9445]<=26'd11119419; ROM3[9445]<=26'd9726757; ROM4[9445]<=26'd23443478;
ROM1[9446]<=26'd1944752; ROM2[9446]<=26'd11108829; ROM3[9446]<=26'd9714050; ROM4[9446]<=26'd23431230;
ROM1[9447]<=26'd1952414; ROM2[9447]<=26'd11107011; ROM3[9447]<=26'd9708180; ROM4[9447]<=26'd23428136;
ROM1[9448]<=26'd1957780; ROM2[9448]<=26'd11104302; ROM3[9448]<=26'd9700670; ROM4[9448]<=26'd23424631;
ROM1[9449]<=26'd1960987; ROM2[9449]<=26'd11108549; ROM3[9449]<=26'd9706210; ROM4[9449]<=26'd23429617;
ROM1[9450]<=26'd1963156; ROM2[9450]<=26'd11117958; ROM3[9450]<=26'd9716363; ROM4[9450]<=26'd23437020;
ROM1[9451]<=26'd1948502; ROM2[9451]<=26'd11111805; ROM3[9451]<=26'd9710433; ROM4[9451]<=26'd23429232;
ROM1[9452]<=26'd1931851; ROM2[9452]<=26'd11102700; ROM3[9452]<=26'd9703672; ROM4[9452]<=26'd23421759;
ROM1[9453]<=26'd1926397; ROM2[9453]<=26'd11101877; ROM3[9453]<=26'd9704074; ROM4[9453]<=26'd23421502;
ROM1[9454]<=26'd1933313; ROM2[9454]<=26'd11105573; ROM3[9454]<=26'd9705744; ROM4[9454]<=26'd23424403;
ROM1[9455]<=26'd1947943; ROM2[9455]<=26'd11109527; ROM3[9455]<=26'd9704201; ROM4[9455]<=26'd23428193;
ROM1[9456]<=26'd1965833; ROM2[9456]<=26'd11115537; ROM3[9456]<=26'd9703346; ROM4[9456]<=26'd23431080;
ROM1[9457]<=26'd1966302; ROM2[9457]<=26'd11116465; ROM3[9457]<=26'd9701139; ROM4[9457]<=26'd23430347;
ROM1[9458]<=26'd1960192; ROM2[9458]<=26'd11116681; ROM3[9458]<=26'd9704153; ROM4[9458]<=26'd23432486;
ROM1[9459]<=26'd1957787; ROM2[9459]<=26'd11120461; ROM3[9459]<=26'd9710889; ROM4[9459]<=26'd23436259;
ROM1[9460]<=26'd1948701; ROM2[9460]<=26'd11114110; ROM3[9460]<=26'd9707436; ROM4[9460]<=26'd23431035;
ROM1[9461]<=26'd1938038; ROM2[9461]<=26'd11107658; ROM3[9461]<=26'd9704854; ROM4[9461]<=26'd23426645;
ROM1[9462]<=26'd1936754; ROM2[9462]<=26'd11106861; ROM3[9462]<=26'd9704221; ROM4[9462]<=26'd23426038;
ROM1[9463]<=26'd1942607; ROM2[9463]<=26'd11106997; ROM3[9463]<=26'd9701660; ROM4[9463]<=26'd23424587;
ROM1[9464]<=26'd1958639; ROM2[9464]<=26'd11113726; ROM3[9464]<=26'd9699855; ROM4[9464]<=26'd23428611;
ROM1[9465]<=26'd1974681; ROM2[9465]<=26'd11125865; ROM3[9465]<=26'd9706981; ROM4[9465]<=26'd23438093;
ROM1[9466]<=26'd1970411; ROM2[9466]<=26'd11126654; ROM3[9466]<=26'd9710799; ROM4[9466]<=26'd23438165;
ROM1[9467]<=26'd1955453; ROM2[9467]<=26'd11116185; ROM3[9467]<=26'd9706492; ROM4[9467]<=26'd23429793;
ROM1[9468]<=26'd1950939; ROM2[9468]<=26'd11116373; ROM3[9468]<=26'd9709609; ROM4[9468]<=26'd23431670;
ROM1[9469]<=26'd1942005; ROM2[9469]<=26'd11114846; ROM3[9469]<=26'd9709593; ROM4[9469]<=26'd23430176;
ROM1[9470]<=26'd1936000; ROM2[9470]<=26'd11111173; ROM3[9470]<=26'd9706574; ROM4[9470]<=26'd23426634;
ROM1[9471]<=26'd1942440; ROM2[9471]<=26'd11112595; ROM3[9471]<=26'd9706202; ROM4[9471]<=26'd23428131;
ROM1[9472]<=26'd1954943; ROM2[9472]<=26'd11113626; ROM3[9472]<=26'd9705446; ROM4[9472]<=26'd23429454;
ROM1[9473]<=26'd1967591; ROM2[9473]<=26'd11118866; ROM3[9473]<=26'd9706985; ROM4[9473]<=26'd23434856;
ROM1[9474]<=26'd1972894; ROM2[9474]<=26'd11125914; ROM3[9474]<=26'd9714715; ROM4[9474]<=26'd23442899;
ROM1[9475]<=26'd1964905; ROM2[9475]<=26'd11122455; ROM3[9475]<=26'd9715958; ROM4[9475]<=26'd23441705;
ROM1[9476]<=26'd1960231; ROM2[9476]<=26'd11122265; ROM3[9476]<=26'd9721107; ROM4[9476]<=26'd23442491;
ROM1[9477]<=26'd1956661; ROM2[9477]<=26'd11121399; ROM3[9477]<=26'd9724527; ROM4[9477]<=26'd23441248;
ROM1[9478]<=26'd1944180; ROM2[9478]<=26'd11113764; ROM3[9478]<=26'd9717906; ROM4[9478]<=26'd23434419;
ROM1[9479]<=26'd1952146; ROM2[9479]<=26'd11120801; ROM3[9479]<=26'd9724405; ROM4[9479]<=26'd23441270;
ROM1[9480]<=26'd1961144; ROM2[9480]<=26'd11118746; ROM3[9480]<=26'd9721048; ROM4[9480]<=26'd23439363;
ROM1[9481]<=26'd1964265; ROM2[9481]<=26'd11109848; ROM3[9481]<=26'd9707569; ROM4[9481]<=26'd23430168;
ROM1[9482]<=26'd1965144; ROM2[9482]<=26'd11108801; ROM3[9482]<=26'd9707308; ROM4[9482]<=26'd23428830;
ROM1[9483]<=26'd1959096; ROM2[9483]<=26'd11109880; ROM3[9483]<=26'd9710341; ROM4[9483]<=26'd23428459;
ROM1[9484]<=26'd1955929; ROM2[9484]<=26'd11114588; ROM3[9484]<=26'd9717021; ROM4[9484]<=26'd23431709;
ROM1[9485]<=26'd1953725; ROM2[9485]<=26'd11116759; ROM3[9485]<=26'd9722067; ROM4[9485]<=26'd23435008;
ROM1[9486]<=26'd1947852; ROM2[9486]<=26'd11115250; ROM3[9486]<=26'd9724158; ROM4[9486]<=26'd23436664;
ROM1[9487]<=26'd1946722; ROM2[9487]<=26'd11114429; ROM3[9487]<=26'd9724535; ROM4[9487]<=26'd23436866;
ROM1[9488]<=26'd1952880; ROM2[9488]<=26'd11115509; ROM3[9488]<=26'd9722054; ROM4[9488]<=26'd23436413;
ROM1[9489]<=26'd1965281; ROM2[9489]<=26'd11116512; ROM3[9489]<=26'd9718417; ROM4[9489]<=26'd23437176;
ROM1[9490]<=26'd1971270; ROM2[9490]<=26'd11117713; ROM3[9490]<=26'd9717749; ROM4[9490]<=26'd23439165;
ROM1[9491]<=26'd1965707; ROM2[9491]<=26'd11116723; ROM3[9491]<=26'd9719967; ROM4[9491]<=26'd23440283;
ROM1[9492]<=26'd1957873; ROM2[9492]<=26'd11116497; ROM3[9492]<=26'd9722402; ROM4[9492]<=26'd23440998;
ROM1[9493]<=26'd1953770; ROM2[9493]<=26'd11117265; ROM3[9493]<=26'd9727638; ROM4[9493]<=26'd23444264;
ROM1[9494]<=26'd1949885; ROM2[9494]<=26'd11116492; ROM3[9494]<=26'd9731600; ROM4[9494]<=26'd23445761;
ROM1[9495]<=26'd1947311; ROM2[9495]<=26'd11114743; ROM3[9495]<=26'd9731175; ROM4[9495]<=26'd23443605;
ROM1[9496]<=26'd1955069; ROM2[9496]<=26'd11116454; ROM3[9496]<=26'd9731328; ROM4[9496]<=26'd23445136;
ROM1[9497]<=26'd1971113; ROM2[9497]<=26'd11120518; ROM3[9497]<=26'd9728098; ROM4[9497]<=26'd23446869;
ROM1[9498]<=26'd1977059; ROM2[9498]<=26'd11118502; ROM3[9498]<=26'd9720368; ROM4[9498]<=26'd23441235;
ROM1[9499]<=26'd1969627; ROM2[9499]<=26'd11113933; ROM3[9499]<=26'd9715692; ROM4[9499]<=26'd23436118;
ROM1[9500]<=26'd1957873; ROM2[9500]<=26'd11111066; ROM3[9500]<=26'd9714197; ROM4[9500]<=26'd23433549;
ROM1[9501]<=26'd1947709; ROM2[9501]<=26'd11107977; ROM3[9501]<=26'd9712760; ROM4[9501]<=26'd23429530;
ROM1[9502]<=26'd1947448; ROM2[9502]<=26'd11113314; ROM3[9502]<=26'd9717961; ROM4[9502]<=26'd23433676;
ROM1[9503]<=26'd1947703; ROM2[9503]<=26'd11118348; ROM3[9503]<=26'd9721344; ROM4[9503]<=26'd23436852;
ROM1[9504]<=26'd1947132; ROM2[9504]<=26'd11114217; ROM3[9504]<=26'd9714949; ROM4[9504]<=26'd23432847;
ROM1[9505]<=26'd1954489; ROM2[9505]<=26'd11112259; ROM3[9505]<=26'd9708478; ROM4[9505]<=26'd23429513;
ROM1[9506]<=26'd1964534; ROM2[9506]<=26'd11111997; ROM3[9506]<=26'd9700807; ROM4[9506]<=26'd23425899;
ROM1[9507]<=26'd1969534; ROM2[9507]<=26'd11117474; ROM3[9507]<=26'd9704656; ROM4[9507]<=26'd23430755;
ROM1[9508]<=26'd1971022; ROM2[9508]<=26'd11123605; ROM3[9508]<=26'd9714862; ROM4[9508]<=26'd23437970;
ROM1[9509]<=26'd1965509; ROM2[9509]<=26'd11123285; ROM3[9509]<=26'd9719006; ROM4[9509]<=26'd23440614;
ROM1[9510]<=26'd1961691; ROM2[9510]<=26'd11125297; ROM3[9510]<=26'd9722368; ROM4[9510]<=26'd23444777;
ROM1[9511]<=26'd1949951; ROM2[9511]<=26'd11116868; ROM3[9511]<=26'd9718918; ROM4[9511]<=26'd23439170;
ROM1[9512]<=26'd1938077; ROM2[9512]<=26'd11105600; ROM3[9512]<=26'd9708483; ROM4[9512]<=26'd23426998;
ROM1[9513]<=26'd1946169; ROM2[9513]<=26'd11108119; ROM3[9513]<=26'd9706006; ROM4[9513]<=26'd23427181;
ROM1[9514]<=26'd1959869; ROM2[9514]<=26'd11110510; ROM3[9514]<=26'd9702522; ROM4[9514]<=26'd23427763;
ROM1[9515]<=26'd1966909; ROM2[9515]<=26'd11113373; ROM3[9515]<=26'd9702317; ROM4[9515]<=26'd23430627;
ROM1[9516]<=26'd1962977; ROM2[9516]<=26'd11112465; ROM3[9516]<=26'd9705034; ROM4[9516]<=26'd23431080;
ROM1[9517]<=26'd1951113; ROM2[9517]<=26'd11106017; ROM3[9517]<=26'd9704125; ROM4[9517]<=26'd23425904;
ROM1[9518]<=26'd1940318; ROM2[9518]<=26'd11101349; ROM3[9518]<=26'd9703741; ROM4[9518]<=26'd23421734;
ROM1[9519]<=26'd1931960; ROM2[9519]<=26'd11097092; ROM3[9519]<=26'd9703910; ROM4[9519]<=26'd23418816;
ROM1[9520]<=26'd1931363; ROM2[9520]<=26'd11098982; ROM3[9520]<=26'd9706673; ROM4[9520]<=26'd23421675;
ROM1[9521]<=26'd1939450; ROM2[9521]<=26'd11103231; ROM3[9521]<=26'd9708600; ROM4[9521]<=26'd23424195;
ROM1[9522]<=26'd1951365; ROM2[9522]<=26'd11104245; ROM3[9522]<=26'd9705438; ROM4[9522]<=26'd23422793;
ROM1[9523]<=26'd1957842; ROM2[9523]<=26'd11102968; ROM3[9523]<=26'd9700400; ROM4[9523]<=26'd23420669;
ROM1[9524]<=26'd1957271; ROM2[9524]<=26'd11104781; ROM3[9524]<=26'd9703055; ROM4[9524]<=26'd23422752;
ROM1[9525]<=26'd1951617; ROM2[9525]<=26'd11106375; ROM3[9525]<=26'd9708088; ROM4[9525]<=26'd23425792;
ROM1[9526]<=26'd1946490; ROM2[9526]<=26'd11105572; ROM3[9526]<=26'd9712409; ROM4[9526]<=26'd23426501;
ROM1[9527]<=26'd1943139; ROM2[9527]<=26'd11107718; ROM3[9527]<=26'd9717131; ROM4[9527]<=26'd23430155;
ROM1[9528]<=26'd1940488; ROM2[9528]<=26'd11111635; ROM3[9528]<=26'd9720670; ROM4[9528]<=26'd23432389;
ROM1[9529]<=26'd1944807; ROM2[9529]<=26'd11112547; ROM3[9529]<=26'd9719180; ROM4[9529]<=26'd23430848;
ROM1[9530]<=26'd1954776; ROM2[9530]<=26'd11113669; ROM3[9530]<=26'd9714729; ROM4[9530]<=26'd23430888;
ROM1[9531]<=26'd1969463; ROM2[9531]<=26'd11117795; ROM3[9531]<=26'd9712971; ROM4[9531]<=26'd23432776;
ROM1[9532]<=26'd1972223; ROM2[9532]<=26'd11115922; ROM3[9532]<=26'd9714226; ROM4[9532]<=26'd23433147;
ROM1[9533]<=26'd1970266; ROM2[9533]<=26'd11119885; ROM3[9533]<=26'd9723657; ROM4[9533]<=26'd23439998;
ROM1[9534]<=26'd1968209; ROM2[9534]<=26'd11123284; ROM3[9534]<=26'd9731582; ROM4[9534]<=26'd23446789;
ROM1[9535]<=26'd1963456; ROM2[9535]<=26'd11121471; ROM3[9535]<=26'd9732979; ROM4[9535]<=26'd23446616;
ROM1[9536]<=26'd1950418; ROM2[9536]<=26'd11112759; ROM3[9536]<=26'd9727945; ROM4[9536]<=26'd23439533;
ROM1[9537]<=26'd1941182; ROM2[9537]<=26'd11102775; ROM3[9537]<=26'd9721789; ROM4[9537]<=26'd23431311;
ROM1[9538]<=26'd1948992; ROM2[9538]<=26'd11104114; ROM3[9538]<=26'd9723992; ROM4[9538]<=26'd23432862;
ROM1[9539]<=26'd1968200; ROM2[9539]<=26'd11111746; ROM3[9539]<=26'd9729538; ROM4[9539]<=26'd23441990;
ROM1[9540]<=26'd1975895; ROM2[9540]<=26'd11113964; ROM3[9540]<=26'd9732566; ROM4[9540]<=26'd23447735;
ROM1[9541]<=26'd1970490; ROM2[9541]<=26'd11112484; ROM3[9541]<=26'd9735682; ROM4[9541]<=26'd23449643;
ROM1[9542]<=26'd1966477; ROM2[9542]<=26'd11113927; ROM3[9542]<=26'd9742645; ROM4[9542]<=26'd23452597;
ROM1[9543]<=26'd1959697; ROM2[9543]<=26'd11110067; ROM3[9543]<=26'd9741654; ROM4[9543]<=26'd23450617;
ROM1[9544]<=26'd1957776; ROM2[9544]<=26'd11113322; ROM3[9544]<=26'd9746691; ROM4[9544]<=26'd23456462;
ROM1[9545]<=26'd1961376; ROM2[9545]<=26'd11120991; ROM3[9545]<=26'd9753833; ROM4[9545]<=26'd23463283;
ROM1[9546]<=26'd1956768; ROM2[9546]<=26'd11112633; ROM3[9546]<=26'd9741125; ROM4[9546]<=26'd23452832;
ROM1[9547]<=26'd1961804; ROM2[9547]<=26'd11107371; ROM3[9547]<=26'd9729240; ROM4[9547]<=26'd23443463;
ROM1[9548]<=26'd1974220; ROM2[9548]<=26'd11112273; ROM3[9548]<=26'd9725886; ROM4[9548]<=26'd23442467;
ROM1[9549]<=26'd1972264; ROM2[9549]<=26'd11113426; ROM3[9549]<=26'd9724291; ROM4[9549]<=26'd23441173;
ROM1[9550]<=26'd1969714; ROM2[9550]<=26'd11118596; ROM3[9550]<=26'd9729488; ROM4[9550]<=26'd23445696;
ROM1[9551]<=26'd1965628; ROM2[9551]<=26'd11121039; ROM3[9551]<=26'd9733322; ROM4[9551]<=26'd23446961;
ROM1[9552]<=26'd1958733; ROM2[9552]<=26'd11120783; ROM3[9552]<=26'd9731152; ROM4[9552]<=26'd23444465;
ROM1[9553]<=26'd1954848; ROM2[9553]<=26'd11119711; ROM3[9553]<=26'd9729358; ROM4[9553]<=26'd23442736;
ROM1[9554]<=26'd1955310; ROM2[9554]<=26'd11119065; ROM3[9554]<=26'd9727245; ROM4[9554]<=26'd23439675;
ROM1[9555]<=26'd1968174; ROM2[9555]<=26'd11123852; ROM3[9555]<=26'd9725810; ROM4[9555]<=26'd23440672;
ROM1[9556]<=26'd1980358; ROM2[9556]<=26'd11125424; ROM3[9556]<=26'd9721821; ROM4[9556]<=26'd23439843;
ROM1[9557]<=26'd1980229; ROM2[9557]<=26'd11125386; ROM3[9557]<=26'd9721237; ROM4[9557]<=26'd23440042;
ROM1[9558]<=26'd1976557; ROM2[9558]<=26'd11126725; ROM3[9558]<=26'd9724981; ROM4[9558]<=26'd23444069;
ROM1[9559]<=26'd1968863; ROM2[9559]<=26'd11124403; ROM3[9559]<=26'd9727033; ROM4[9559]<=26'd23443632;
ROM1[9560]<=26'd1962380; ROM2[9560]<=26'd11122661; ROM3[9560]<=26'd9727853; ROM4[9560]<=26'd23443205;
ROM1[9561]<=26'd1953719; ROM2[9561]<=26'd11119899; ROM3[9561]<=26'd9727451; ROM4[9561]<=26'd23440305;
ROM1[9562]<=26'd1951633; ROM2[9562]<=26'd11116667; ROM3[9562]<=26'd9724928; ROM4[9562]<=26'd23437659;
ROM1[9563]<=26'd1958572; ROM2[9563]<=26'd11119500; ROM3[9563]<=26'd9721066; ROM4[9563]<=26'd23438800;
ROM1[9564]<=26'd1971902; ROM2[9564]<=26'd11122994; ROM3[9564]<=26'd9718678; ROM4[9564]<=26'd23440300;
ROM1[9565]<=26'd1977631; ROM2[9565]<=26'd11121600; ROM3[9565]<=26'd9716790; ROM4[9565]<=26'd23441485;
ROM1[9566]<=26'd1973016; ROM2[9566]<=26'd11121458; ROM3[9566]<=26'd9719004; ROM4[9566]<=26'd23443229;
ROM1[9567]<=26'd1967947; ROM2[9567]<=26'd11124593; ROM3[9567]<=26'd9723542; ROM4[9567]<=26'd23447364;
ROM1[9568]<=26'd1966057; ROM2[9568]<=26'd11129595; ROM3[9568]<=26'd9729801; ROM4[9568]<=26'd23452461;
ROM1[9569]<=26'd1959839; ROM2[9569]<=26'd11129771; ROM3[9569]<=26'd9732122; ROM4[9569]<=26'd23452416;
ROM1[9570]<=26'd1959053; ROM2[9570]<=26'd11130602; ROM3[9570]<=26'd9733738; ROM4[9570]<=26'd23453336;
ROM1[9571]<=26'd1963343; ROM2[9571]<=26'd11128765; ROM3[9571]<=26'd9731613; ROM4[9571]<=26'd23451117;
ROM1[9572]<=26'd1966145; ROM2[9572]<=26'd11120357; ROM3[9572]<=26'd9718388; ROM4[9572]<=26'd23441641;
ROM1[9573]<=26'd1972416; ROM2[9573]<=26'd11120141; ROM3[9573]<=26'd9710751; ROM4[9573]<=26'd23438754;
ROM1[9574]<=26'd1967104; ROM2[9574]<=26'd11118074; ROM3[9574]<=26'd9708219; ROM4[9574]<=26'd23434769;
ROM1[9575]<=26'd1951443; ROM2[9575]<=26'd11108387; ROM3[9575]<=26'd9702930; ROM4[9575]<=26'd23425452;
ROM1[9576]<=26'd1942445; ROM2[9576]<=26'd11102456; ROM3[9576]<=26'd9703999; ROM4[9576]<=26'd23421321;
ROM1[9577]<=26'd1938459; ROM2[9577]<=26'd11102153; ROM3[9577]<=26'd9708124; ROM4[9577]<=26'd23420928;
ROM1[9578]<=26'd1935133; ROM2[9578]<=26'd11103471; ROM3[9578]<=26'd9709335; ROM4[9578]<=26'd23420886;
ROM1[9579]<=26'd1941484; ROM2[9579]<=26'd11108482; ROM3[9579]<=26'd9712356; ROM4[9579]<=26'd23424250;
ROM1[9580]<=26'd1953629; ROM2[9580]<=26'd11113091; ROM3[9580]<=26'd9711061; ROM4[9580]<=26'd23425081;
ROM1[9581]<=26'd1964543; ROM2[9581]<=26'd11112463; ROM3[9581]<=26'd9705674; ROM4[9581]<=26'd23423573;
ROM1[9582]<=26'd1968076; ROM2[9582]<=26'd11114149; ROM3[9582]<=26'd9709872; ROM4[9582]<=26'd23426467;
ROM1[9583]<=26'd1966497; ROM2[9583]<=26'd11120939; ROM3[9583]<=26'd9718309; ROM4[9583]<=26'd23432078;
ROM1[9584]<=26'd1949762; ROM2[9584]<=26'd11109750; ROM3[9584]<=26'd9712571; ROM4[9584]<=26'd23423336;
ROM1[9585]<=26'd1936404; ROM2[9585]<=26'd11099050; ROM3[9585]<=26'd9707016; ROM4[9585]<=26'd23415027;
ROM1[9586]<=26'd1928906; ROM2[9586]<=26'd11096284; ROM3[9586]<=26'd9705952; ROM4[9586]<=26'd23413151;
ROM1[9587]<=26'd1927206; ROM2[9587]<=26'd11092425; ROM3[9587]<=26'd9704477; ROM4[9587]<=26'd23410483;
ROM1[9588]<=26'd1942184; ROM2[9588]<=26'd11099399; ROM3[9588]<=26'd9710211; ROM4[9588]<=26'd23417329;
ROM1[9589]<=26'd1959229; ROM2[9589]<=26'd11105276; ROM3[9589]<=26'd9710021; ROM4[9589]<=26'd23423403;
ROM1[9590]<=26'd1962252; ROM2[9590]<=26'd11103801; ROM3[9590]<=26'd9707183; ROM4[9590]<=26'd23423171;
ROM1[9591]<=26'd1955940; ROM2[9591]<=26'd11100299; ROM3[9591]<=26'd9710595; ROM4[9591]<=26'd23425922;
ROM1[9592]<=26'd1953994; ROM2[9592]<=26'd11104063; ROM3[9592]<=26'd9717697; ROM4[9592]<=26'd23432507;
ROM1[9593]<=26'd1953440; ROM2[9593]<=26'd11109302; ROM3[9593]<=26'd9726849; ROM4[9593]<=26'd23439123;
ROM1[9594]<=26'd1949817; ROM2[9594]<=26'd11110750; ROM3[9594]<=26'd9735318; ROM4[9594]<=26'd23443997;
ROM1[9595]<=26'd1949654; ROM2[9595]<=26'd11110831; ROM3[9595]<=26'd9738556; ROM4[9595]<=26'd23446515;
ROM1[9596]<=26'd1955620; ROM2[9596]<=26'd11110668; ROM3[9596]<=26'd9739238; ROM4[9596]<=26'd23448554;
ROM1[9597]<=26'd1968286; ROM2[9597]<=26'd11112314; ROM3[9597]<=26'd9737875; ROM4[9597]<=26'd23451047;
ROM1[9598]<=26'd1978714; ROM2[9598]<=26'd11114063; ROM3[9598]<=26'd9736856; ROM4[9598]<=26'd23453707;
ROM1[9599]<=26'd1978351; ROM2[9599]<=26'd11115914; ROM3[9599]<=26'd9740348; ROM4[9599]<=26'd23456594;
ROM1[9600]<=26'd1973918; ROM2[9600]<=26'd11118644; ROM3[9600]<=26'd9747064; ROM4[9600]<=26'd23460807;
ROM1[9601]<=26'd1970238; ROM2[9601]<=26'd11121173; ROM3[9601]<=26'd9753413; ROM4[9601]<=26'd23462224;
ROM1[9602]<=26'd1966405; ROM2[9602]<=26'd11120510; ROM3[9602]<=26'd9756275; ROM4[9602]<=26'd23463409;
ROM1[9603]<=26'd1959861; ROM2[9603]<=26'd11118876; ROM3[9603]<=26'd9755261; ROM4[9603]<=26'd23459494;
ROM1[9604]<=26'd1963589; ROM2[9604]<=26'd11123686; ROM3[9604]<=26'd9756955; ROM4[9604]<=26'd23460418;
ROM1[9605]<=26'd1971085; ROM2[9605]<=26'd11120452; ROM3[9605]<=26'd9747035; ROM4[9605]<=26'd23455465;
ROM1[9606]<=26'd1975138; ROM2[9606]<=26'd11114399; ROM3[9606]<=26'd9730977; ROM4[9606]<=26'd23444384;
ROM1[9607]<=26'd1976076; ROM2[9607]<=26'd11114290; ROM3[9607]<=26'd9726923; ROM4[9607]<=26'd23443043;
ROM1[9608]<=26'd1969528; ROM2[9608]<=26'd11112867; ROM3[9608]<=26'd9726611; ROM4[9608]<=26'd23440846;
ROM1[9609]<=26'd1967556; ROM2[9609]<=26'd11117667; ROM3[9609]<=26'd9732838; ROM4[9609]<=26'd23444216;
ROM1[9610]<=26'd1972043; ROM2[9610]<=26'd11125568; ROM3[9610]<=26'd9741648; ROM4[9610]<=26'd23449608;
ROM1[9611]<=26'd1963299; ROM2[9611]<=26'd11120722; ROM3[9611]<=26'd9739217; ROM4[9611]<=26'd23443165;
ROM1[9612]<=26'd1954279; ROM2[9612]<=26'd11111213; ROM3[9612]<=26'd9727909; ROM4[9612]<=26'd23433431;
ROM1[9613]<=26'd1959058; ROM2[9613]<=26'd11109023; ROM3[9613]<=26'd9718972; ROM4[9613]<=26'd23428235;
ROM1[9614]<=26'd1968833; ROM2[9614]<=26'd11107075; ROM3[9614]<=26'd9710250; ROM4[9614]<=26'd23423607;
ROM1[9615]<=26'd1974922; ROM2[9615]<=26'd11107572; ROM3[9615]<=26'd9706566; ROM4[9615]<=26'd23423928;
ROM1[9616]<=26'd1973929; ROM2[9616]<=26'd11110443; ROM3[9616]<=26'd9709782; ROM4[9616]<=26'd23426058;
ROM1[9617]<=26'd1969699; ROM2[9617]<=26'd11113618; ROM3[9617]<=26'd9719407; ROM4[9617]<=26'd23430040;
ROM1[9618]<=26'd1959750; ROM2[9618]<=26'd11110381; ROM3[9618]<=26'd9717355; ROM4[9618]<=26'd23426026;
ROM1[9619]<=26'd1949618; ROM2[9619]<=26'd11107567; ROM3[9619]<=26'd9715368; ROM4[9619]<=26'd23422538;
ROM1[9620]<=26'd1949386; ROM2[9620]<=26'd11111073; ROM3[9620]<=26'd9718381; ROM4[9620]<=26'd23425325;
ROM1[9621]<=26'd1950171; ROM2[9621]<=26'd11108314; ROM3[9621]<=26'd9709085; ROM4[9621]<=26'd23418484;
ROM1[9622]<=26'd1958545; ROM2[9622]<=26'd11109139; ROM3[9622]<=26'd9700993; ROM4[9622]<=26'd23416347;
ROM1[9623]<=26'd1969006; ROM2[9623]<=26'd11115743; ROM3[9623]<=26'd9698694; ROM4[9623]<=26'd23419919;
ROM1[9624]<=26'd1967163; ROM2[9624]<=26'd11115903; ROM3[9624]<=26'd9699460; ROM4[9624]<=26'd23419931;
ROM1[9625]<=26'd1956101; ROM2[9625]<=26'd11110838; ROM3[9625]<=26'd9700025; ROM4[9625]<=26'd23418763;
ROM1[9626]<=26'd1950338; ROM2[9626]<=26'd11112320; ROM3[9626]<=26'd9706312; ROM4[9626]<=26'd23423268;
ROM1[9627]<=26'd1948589; ROM2[9627]<=26'd11114024; ROM3[9627]<=26'd9714219; ROM4[9627]<=26'd23427576;
ROM1[9628]<=26'd1943709; ROM2[9628]<=26'd11111879; ROM3[9628]<=26'd9714576; ROM4[9628]<=26'd23427198;
ROM1[9629]<=26'd1946297; ROM2[9629]<=26'd11113564; ROM3[9629]<=26'd9715483; ROM4[9629]<=26'd23429159;
ROM1[9630]<=26'd1959077; ROM2[9630]<=26'd11116438; ROM3[9630]<=26'd9715796; ROM4[9630]<=26'd23429979;
ROM1[9631]<=26'd1973340; ROM2[9631]<=26'd11117976; ROM3[9631]<=26'd9713938; ROM4[9631]<=26'd23432258;
ROM1[9632]<=26'd1975114; ROM2[9632]<=26'd11118318; ROM3[9632]<=26'd9715781; ROM4[9632]<=26'd23434804;
ROM1[9633]<=26'd1971094; ROM2[9633]<=26'd11119371; ROM3[9633]<=26'd9723371; ROM4[9633]<=26'd23438421;
ROM1[9634]<=26'd1966274; ROM2[9634]<=26'd11116527; ROM3[9634]<=26'd9730703; ROM4[9634]<=26'd23442365;
ROM1[9635]<=26'd1961495; ROM2[9635]<=26'd11113368; ROM3[9635]<=26'd9733498; ROM4[9635]<=26'd23442595;
ROM1[9636]<=26'd1956586; ROM2[9636]<=26'd11112385; ROM3[9636]<=26'd9738553; ROM4[9636]<=26'd23443490;
ROM1[9637]<=26'd1958703; ROM2[9637]<=26'd11112396; ROM3[9637]<=26'd9740223; ROM4[9637]<=26'd23445561;
ROM1[9638]<=26'd1969960; ROM2[9638]<=26'd11116175; ROM3[9638]<=26'd9740263; ROM4[9638]<=26'd23448022;
ROM1[9639]<=26'd1984150; ROM2[9639]<=26'd11118297; ROM3[9639]<=26'd9736947; ROM4[9639]<=26'd23447819;
ROM1[9640]<=26'd1990774; ROM2[9640]<=26'd11117473; ROM3[9640]<=26'd9736879; ROM4[9640]<=26'd23448447;
ROM1[9641]<=26'd1991618; ROM2[9641]<=26'd11120207; ROM3[9641]<=26'd9744537; ROM4[9641]<=26'd23454264;
ROM1[9642]<=26'd1977416; ROM2[9642]<=26'd11113382; ROM3[9642]<=26'd9740940; ROM4[9642]<=26'd23448205;
ROM1[9643]<=26'd1966184; ROM2[9643]<=26'd11106170; ROM3[9643]<=26'd9736881; ROM4[9643]<=26'd23440423;
ROM1[9644]<=26'd1967900; ROM2[9644]<=26'd11112355; ROM3[9644]<=26'd9746143; ROM4[9644]<=26'd23447332;
ROM1[9645]<=26'd1962547; ROM2[9645]<=26'd11109476; ROM3[9645]<=26'd9744938; ROM4[9645]<=26'd23444094;
ROM1[9646]<=26'd1964848; ROM2[9646]<=26'd11105918; ROM3[9646]<=26'd9739997; ROM4[9646]<=26'd23441371;
ROM1[9647]<=26'd1974020; ROM2[9647]<=26'd11103929; ROM3[9647]<=26'd9733717; ROM4[9647]<=26'd23440155;
ROM1[9648]<=26'd1972253; ROM2[9648]<=26'd11094656; ROM3[9648]<=26'd9719314; ROM4[9648]<=26'd23429101;
ROM1[9649]<=26'd1965483; ROM2[9649]<=26'd11092038; ROM3[9649]<=26'd9714948; ROM4[9649]<=26'd23426218;
ROM1[9650]<=26'd1961617; ROM2[9650]<=26'd11096066; ROM3[9650]<=26'd9721433; ROM4[9650]<=26'd23430441;
ROM1[9651]<=26'd1959678; ROM2[9651]<=26'd11100704; ROM3[9651]<=26'd9727533; ROM4[9651]<=26'd23435009;
ROM1[9652]<=26'd1957537; ROM2[9652]<=26'd11103727; ROM3[9652]<=26'd9730907; ROM4[9652]<=26'd23437163;
ROM1[9653]<=26'd1954277; ROM2[9653]<=26'd11104502; ROM3[9653]<=26'd9732957; ROM4[9653]<=26'd23436654;
ROM1[9654]<=26'd1962973; ROM2[9654]<=26'd11109712; ROM3[9654]<=26'd9737428; ROM4[9654]<=26'd23441502;
ROM1[9655]<=26'd1979531; ROM2[9655]<=26'd11116728; ROM3[9655]<=26'd9739862; ROM4[9655]<=26'd23447342;
ROM1[9656]<=26'd1984357; ROM2[9656]<=26'd11111645; ROM3[9656]<=26'd9726886; ROM4[9656]<=26'd23440659;
ROM1[9657]<=26'd1978172; ROM2[9657]<=26'd11103610; ROM3[9657]<=26'd9714709; ROM4[9657]<=26'd23431017;
ROM1[9658]<=26'd1968009; ROM2[9658]<=26'd11100189; ROM3[9658]<=26'd9709269; ROM4[9658]<=26'd23424861;
ROM1[9659]<=26'd1958701; ROM2[9659]<=26'd11098490; ROM3[9659]<=26'd9708799; ROM4[9659]<=26'd23422616;
ROM1[9660]<=26'd1954519; ROM2[9660]<=26'd11099523; ROM3[9660]<=26'd9712690; ROM4[9660]<=26'd23424795;
ROM1[9661]<=26'd1949218; ROM2[9661]<=26'd11098873; ROM3[9661]<=26'd9714297; ROM4[9661]<=26'd23425432;
ROM1[9662]<=26'd1948610; ROM2[9662]<=26'd11097482; ROM3[9662]<=26'd9711250; ROM4[9662]<=26'd23423139;
ROM1[9663]<=26'd1957098; ROM2[9663]<=26'd11100995; ROM3[9663]<=26'd9706334; ROM4[9663]<=26'd23421826;
ROM1[9664]<=26'd1971923; ROM2[9664]<=26'd11106774; ROM3[9664]<=26'd9701887; ROM4[9664]<=26'd23422624;
ROM1[9665]<=26'd1980805; ROM2[9665]<=26'd11112943; ROM3[9665]<=26'd9702636; ROM4[9665]<=26'd23426685;
ROM1[9666]<=26'd1977914; ROM2[9666]<=26'd11115674; ROM3[9666]<=26'd9706036; ROM4[9666]<=26'd23429995;
ROM1[9667]<=26'd1972074; ROM2[9667]<=26'd11118357; ROM3[9667]<=26'd9712865; ROM4[9667]<=26'd23433243;
ROM1[9668]<=26'd1974757; ROM2[9668]<=26'd11126854; ROM3[9668]<=26'd9723340; ROM4[9668]<=26'd23440995;
ROM1[9669]<=26'd1966939; ROM2[9669]<=26'd11125370; ROM3[9669]<=26'd9724570; ROM4[9669]<=26'd23438878;
ROM1[9670]<=26'd1956267; ROM2[9670]<=26'd11116972; ROM3[9670]<=26'd9717615; ROM4[9670]<=26'd23431144;
ROM1[9671]<=26'd1955506; ROM2[9671]<=26'd11109741; ROM3[9671]<=26'd9710773; ROM4[9671]<=26'd23424715;
ROM1[9672]<=26'd1964060; ROM2[9672]<=26'd11107301; ROM3[9672]<=26'd9704620; ROM4[9672]<=26'd23421594;
ROM1[9673]<=26'd1977666; ROM2[9673]<=26'd11112042; ROM3[9673]<=26'd9704070; ROM4[9673]<=26'd23425904;
ROM1[9674]<=26'd1978001; ROM2[9674]<=26'd11113057; ROM3[9674]<=26'd9708925; ROM4[9674]<=26'd23428645;
ROM1[9675]<=26'd1973537; ROM2[9675]<=26'd11114138; ROM3[9675]<=26'd9716950; ROM4[9675]<=26'd23431935;
ROM1[9676]<=26'd1964069; ROM2[9676]<=26'd11109903; ROM3[9676]<=26'd9719149; ROM4[9676]<=26'd23429773;
ROM1[9677]<=26'd1953697; ROM2[9677]<=26'd11104620; ROM3[9677]<=26'd9719470; ROM4[9677]<=26'd23425845;
ROM1[9678]<=26'd1951600; ROM2[9678]<=26'd11108087; ROM3[9678]<=26'd9724992; ROM4[9678]<=26'd23428776;
ROM1[9679]<=26'd1955684; ROM2[9679]<=26'd11109713; ROM3[9679]<=26'd9725843; ROM4[9679]<=26'd23430675;
ROM1[9680]<=26'd1969683; ROM2[9680]<=26'd11112956; ROM3[9680]<=26'd9726203; ROM4[9680]<=26'd23434890;
ROM1[9681]<=26'd1984983; ROM2[9681]<=26'd11115943; ROM3[9681]<=26'd9724843; ROM4[9681]<=26'd23438653;
ROM1[9682]<=26'd1986866; ROM2[9682]<=26'd11115624; ROM3[9682]<=26'd9726378; ROM4[9682]<=26'd23440616;
ROM1[9683]<=26'd1985527; ROM2[9683]<=26'd11119446; ROM3[9683]<=26'd9735555; ROM4[9683]<=26'd23447872;
ROM1[9684]<=26'd1984784; ROM2[9684]<=26'd11125861; ROM3[9684]<=26'd9744597; ROM4[9684]<=26'd23455616;
ROM1[9685]<=26'd1972538; ROM2[9685]<=26'd11119913; ROM3[9685]<=26'd9742728; ROM4[9685]<=26'd23450821;
ROM1[9686]<=26'd1956619; ROM2[9686]<=26'd11108090; ROM3[9686]<=26'd9734551; ROM4[9686]<=26'd23441247;
ROM1[9687]<=26'd1955133; ROM2[9687]<=26'd11106028; ROM3[9687]<=26'd9731655; ROM4[9687]<=26'd23439127;
ROM1[9688]<=26'd1960800; ROM2[9688]<=26'd11104315; ROM3[9688]<=26'd9727505; ROM4[9688]<=26'd23436718;
ROM1[9689]<=26'd1978407; ROM2[9689]<=26'd11109538; ROM3[9689]<=26'd9727046; ROM4[9689]<=26'd23441013;
ROM1[9690]<=26'd1991505; ROM2[9690]<=26'd11117323; ROM3[9690]<=26'd9732328; ROM4[9690]<=26'd23447210;
ROM1[9691]<=26'd1990191; ROM2[9691]<=26'd11120341; ROM3[9691]<=26'd9735651; ROM4[9691]<=26'd23449909;
ROM1[9692]<=26'd1984156; ROM2[9692]<=26'd11121955; ROM3[9692]<=26'd9740778; ROM4[9692]<=26'd23453214;
ROM1[9693]<=26'd1969914; ROM2[9693]<=26'd11112505; ROM3[9693]<=26'd9737141; ROM4[9693]<=26'd23443640;
ROM1[9694]<=26'd1950918; ROM2[9694]<=26'd11096741; ROM3[9694]<=26'd9724156; ROM4[9694]<=26'd23429113;
ROM1[9695]<=26'd1939403; ROM2[9695]<=26'd11086017; ROM3[9695]<=26'd9716402; ROM4[9695]<=26'd23420122;
ROM1[9696]<=26'd1940799; ROM2[9696]<=26'd11083107; ROM3[9696]<=26'd9711306; ROM4[9696]<=26'd23415800;
ROM1[9697]<=26'd1961313; ROM2[9697]<=26'd11091455; ROM3[9697]<=26'd9712850; ROM4[9697]<=26'd23424149;
ROM1[9698]<=26'd1979869; ROM2[9698]<=26'd11102284; ROM3[9698]<=26'd9720075; ROM4[9698]<=26'd23433467;
ROM1[9699]<=26'd1977696; ROM2[9699]<=26'd11104003; ROM3[9699]<=26'd9721226; ROM4[9699]<=26'd23433587;
ROM1[9700]<=26'd1967577; ROM2[9700]<=26'd11098969; ROM3[9700]<=26'd9716601; ROM4[9700]<=26'd23428800;
ROM1[9701]<=26'd1970032; ROM2[9701]<=26'd11108191; ROM3[9701]<=26'd9725718; ROM4[9701]<=26'd23437413;
ROM1[9702]<=26'd1969914; ROM2[9702]<=26'd11115199; ROM3[9702]<=26'd9735841; ROM4[9702]<=26'd23444400;
ROM1[9703]<=26'd1958350; ROM2[9703]<=26'd11108424; ROM3[9703]<=26'd9731969; ROM4[9703]<=26'd23438403;
ROM1[9704]<=26'd1957699; ROM2[9704]<=26'd11105038; ROM3[9704]<=26'd9726475; ROM4[9704]<=26'd23434378;
ROM1[9705]<=26'd1964906; ROM2[9705]<=26'd11101785; ROM3[9705]<=26'd9718491; ROM4[9705]<=26'd23429202;
ROM1[9706]<=26'd1975634; ROM2[9706]<=26'd11102755; ROM3[9706]<=26'd9712373; ROM4[9706]<=26'd23427461;
ROM1[9707]<=26'd1977707; ROM2[9707]<=26'd11106758; ROM3[9707]<=26'd9713315; ROM4[9707]<=26'd23429835;
ROM1[9708]<=26'd1972567; ROM2[9708]<=26'd11107699; ROM3[9708]<=26'd9718615; ROM4[9708]<=26'd23431803;
ROM1[9709]<=26'd1966595; ROM2[9709]<=26'd11109238; ROM3[9709]<=26'd9723100; ROM4[9709]<=26'd23433233;
ROM1[9710]<=26'd1964051; ROM2[9710]<=26'd11112615; ROM3[9710]<=26'd9727813; ROM4[9710]<=26'd23437528;
ROM1[9711]<=26'd1961292; ROM2[9711]<=26'd11112215; ROM3[9711]<=26'd9731130; ROM4[9711]<=26'd23438878;
ROM1[9712]<=26'd1964138; ROM2[9712]<=26'd11117414; ROM3[9712]<=26'd9736796; ROM4[9712]<=26'd23442872;
ROM1[9713]<=26'd1974727; ROM2[9713]<=26'd11124223; ROM3[9713]<=26'd9739720; ROM4[9713]<=26'd23448796;
ROM1[9714]<=26'd1982593; ROM2[9714]<=26'd11121979; ROM3[9714]<=26'd9728180; ROM4[9714]<=26'd23443649;
ROM1[9715]<=26'd1982989; ROM2[9715]<=26'd11119917; ROM3[9715]<=26'd9720938; ROM4[9715]<=26'd23440028;
ROM1[9716]<=26'd1976340; ROM2[9716]<=26'd11117209; ROM3[9716]<=26'd9721508; ROM4[9716]<=26'd23437560;
ROM1[9717]<=26'd1964795; ROM2[9717]<=26'd11111923; ROM3[9717]<=26'd9720900; ROM4[9717]<=26'd23432669;
ROM1[9718]<=26'd1960272; ROM2[9718]<=26'd11112101; ROM3[9718]<=26'd9724350; ROM4[9718]<=26'd23435754;
ROM1[9719]<=26'd1957923; ROM2[9719]<=26'd11114618; ROM3[9719]<=26'd9729550; ROM4[9719]<=26'd23439691;
ROM1[9720]<=26'd1958050; ROM2[9720]<=26'd11116531; ROM3[9720]<=26'd9728698; ROM4[9720]<=26'd23441208;
ROM1[9721]<=26'd1965060; ROM2[9721]<=26'd11117088; ROM3[9721]<=26'd9726334; ROM4[9721]<=26'd23441117;
ROM1[9722]<=26'd1980788; ROM2[9722]<=26'd11118785; ROM3[9722]<=26'd9725722; ROM4[9722]<=26'd23442440;
ROM1[9723]<=26'd1983656; ROM2[9723]<=26'd11112147; ROM3[9723]<=26'd9715705; ROM4[9723]<=26'd23436203;
ROM1[9724]<=26'd1971966; ROM2[9724]<=26'd11101426; ROM3[9724]<=26'd9708970; ROM4[9724]<=26'd23428873;
ROM1[9725]<=26'd1962840; ROM2[9725]<=26'd11100283; ROM3[9725]<=26'd9710540; ROM4[9725]<=26'd23428670;
ROM1[9726]<=26'd1958029; ROM2[9726]<=26'd11101965; ROM3[9726]<=26'd9714978; ROM4[9726]<=26'd23429016;
ROM1[9727]<=26'd1965130; ROM2[9727]<=26'd11112457; ROM3[9727]<=26'd9729540; ROM4[9727]<=26'd23441326;
ROM1[9728]<=26'd1971169; ROM2[9728]<=26'd11121402; ROM3[9728]<=26'd9738729; ROM4[9728]<=26'd23451493;
ROM1[9729]<=26'd1969023; ROM2[9729]<=26'd11112854; ROM3[9729]<=26'd9730455; ROM4[9729]<=26'd23443713;
ROM1[9730]<=26'd1976382; ROM2[9730]<=26'd11110856; ROM3[9730]<=26'd9723757; ROM4[9730]<=26'd23440522;
ROM1[9731]<=26'd1991297; ROM2[9731]<=26'd11117824; ROM3[9731]<=26'd9723068; ROM4[9731]<=26'd23445383;
ROM1[9732]<=26'd1988280; ROM2[9732]<=26'd11115533; ROM3[9732]<=26'd9721020; ROM4[9732]<=26'd23442211;
ROM1[9733]<=26'd1977887; ROM2[9733]<=26'd11112426; ROM3[9733]<=26'd9719789; ROM4[9733]<=26'd23438952;
ROM1[9734]<=26'd1968903; ROM2[9734]<=26'd11111639; ROM3[9734]<=26'd9720479; ROM4[9734]<=26'd23438429;
ROM1[9735]<=26'd1962471; ROM2[9735]<=26'd11112149; ROM3[9735]<=26'd9721344; ROM4[9735]<=26'd23435717;
ROM1[9736]<=26'd1957505; ROM2[9736]<=26'd11111485; ROM3[9736]<=26'd9719973; ROM4[9736]<=26'd23435096;
ROM1[9737]<=26'd1961234; ROM2[9737]<=26'd11114071; ROM3[9737]<=26'd9722556; ROM4[9737]<=26'd23438029;
ROM1[9738]<=26'd1970930; ROM2[9738]<=26'd11117197; ROM3[9738]<=26'd9722045; ROM4[9738]<=26'd23439172;
ROM1[9739]<=26'd1981853; ROM2[9739]<=26'd11117774; ROM3[9739]<=26'd9715807; ROM4[9739]<=26'd23437579;
ROM1[9740]<=26'd1987753; ROM2[9740]<=26'd11119466; ROM3[9740]<=26'd9714840; ROM4[9740]<=26'd23437831;
ROM1[9741]<=26'd1982234; ROM2[9741]<=26'd11120719; ROM3[9741]<=26'd9718230; ROM4[9741]<=26'd23440087;
ROM1[9742]<=26'd1976385; ROM2[9742]<=26'd11121197; ROM3[9742]<=26'd9723921; ROM4[9742]<=26'd23440995;
ROM1[9743]<=26'd1975525; ROM2[9743]<=26'd11121536; ROM3[9743]<=26'd9730050; ROM4[9743]<=26'd23444520;
ROM1[9744]<=26'd1966073; ROM2[9744]<=26'd11117815; ROM3[9744]<=26'd9729819; ROM4[9744]<=26'd23443035;
ROM1[9745]<=26'd1958423; ROM2[9745]<=26'd11112969; ROM3[9745]<=26'd9725934; ROM4[9745]<=26'd23439308;
ROM1[9746]<=26'd1961136; ROM2[9746]<=26'd11110370; ROM3[9746]<=26'd9721425; ROM4[9746]<=26'd23438003;
ROM1[9747]<=26'd1970161; ROM2[9747]<=26'd11109359; ROM3[9747]<=26'd9714108; ROM4[9747]<=26'd23434052;
ROM1[9748]<=26'd1978898; ROM2[9748]<=26'd11112049; ROM3[9748]<=26'd9714432; ROM4[9748]<=26'd23435801;
ROM1[9749]<=26'd1976824; ROM2[9749]<=26'd11114005; ROM3[9749]<=26'd9718596; ROM4[9749]<=26'd23438066;
ROM1[9750]<=26'd1969490; ROM2[9750]<=26'd11113144; ROM3[9750]<=26'd9722044; ROM4[9750]<=26'd23438027;
ROM1[9751]<=26'd1963261; ROM2[9751]<=26'd11108948; ROM3[9751]<=26'd9723565; ROM4[9751]<=26'd23437059;
ROM1[9752]<=26'd1959722; ROM2[9752]<=26'd11108590; ROM3[9752]<=26'd9725574; ROM4[9752]<=26'd23438044;
ROM1[9753]<=26'd1958218; ROM2[9753]<=26'd11110776; ROM3[9753]<=26'd9730710; ROM4[9753]<=26'd23440803;
ROM1[9754]<=26'd1959344; ROM2[9754]<=26'd11111476; ROM3[9754]<=26'd9732666; ROM4[9754]<=26'd23441520;
ROM1[9755]<=26'd1965192; ROM2[9755]<=26'd11111005; ROM3[9755]<=26'd9726168; ROM4[9755]<=26'd23439630;
ROM1[9756]<=26'd1975694; ROM2[9756]<=26'd11111650; ROM3[9756]<=26'd9719013; ROM4[9756]<=26'd23437332;
ROM1[9757]<=26'd1980764; ROM2[9757]<=26'd11113513; ROM3[9757]<=26'd9719507; ROM4[9757]<=26'd23438405;
ROM1[9758]<=26'd1977654; ROM2[9758]<=26'd11115241; ROM3[9758]<=26'd9722078; ROM4[9758]<=26'd23440606;
ROM1[9759]<=26'd1967576; ROM2[9759]<=26'd11112187; ROM3[9759]<=26'd9725409; ROM4[9759]<=26'd23439942;
ROM1[9760]<=26'd1961717; ROM2[9760]<=26'd11111585; ROM3[9760]<=26'd9728930; ROM4[9760]<=26'd23440563;
ROM1[9761]<=26'd1963854; ROM2[9761]<=26'd11118670; ROM3[9761]<=26'd9736687; ROM4[9761]<=26'd23447699;
ROM1[9762]<=26'd1963823; ROM2[9762]<=26'd11117450; ROM3[9762]<=26'd9733481; ROM4[9762]<=26'd23446803;
ROM1[9763]<=26'd1962593; ROM2[9763]<=26'd11109049; ROM3[9763]<=26'd9717871; ROM4[9763]<=26'd23434560;
ROM1[9764]<=26'd1977507; ROM2[9764]<=26'd11111967; ROM3[9764]<=26'd9714270; ROM4[9764]<=26'd23434667;
ROM1[9765]<=26'd1984484; ROM2[9765]<=26'd11114839; ROM3[9765]<=26'd9713209; ROM4[9765]<=26'd23436466;
ROM1[9766]<=26'd1981000; ROM2[9766]<=26'd11117258; ROM3[9766]<=26'd9715397; ROM4[9766]<=26'd23436471;
ROM1[9767]<=26'd1980797; ROM2[9767]<=26'd11123638; ROM3[9767]<=26'd9724308; ROM4[9767]<=26'd23443132;
ROM1[9768]<=26'd1978214; ROM2[9768]<=26'd11124879; ROM3[9768]<=26'd9727172; ROM4[9768]<=26'd23445016;
ROM1[9769]<=26'd1966760; ROM2[9769]<=26'd11120423; ROM3[9769]<=26'd9723610; ROM4[9769]<=26'd23439221;
ROM1[9770]<=26'd1963572; ROM2[9770]<=26'd11119991; ROM3[9770]<=26'd9723099; ROM4[9770]<=26'd23437253;
ROM1[9771]<=26'd1972816; ROM2[9771]<=26'd11123733; ROM3[9771]<=26'd9722926; ROM4[9771]<=26'd23439043;
ROM1[9772]<=26'd1984937; ROM2[9772]<=26'd11124991; ROM3[9772]<=26'd9716915; ROM4[9772]<=26'd23437354;
ROM1[9773]<=26'd1994668; ROM2[9773]<=26'd11125339; ROM3[9773]<=26'd9713775; ROM4[9773]<=26'd23437941;
ROM1[9774]<=26'd1998598; ROM2[9774]<=26'd11132418; ROM3[9774]<=26'd9722595; ROM4[9774]<=26'd23446874;
ROM1[9775]<=26'd2002489; ROM2[9775]<=26'd11144664; ROM3[9775]<=26'd9737520; ROM4[9775]<=26'd23459963;
ROM1[9776]<=26'd1988004; ROM2[9776]<=26'd11135757; ROM3[9776]<=26'd9732121; ROM4[9776]<=26'd23451365;
ROM1[9777]<=26'd1971513; ROM2[9777]<=26'd11123358; ROM3[9777]<=26'd9724307; ROM4[9777]<=26'd23439181;
ROM1[9778]<=26'd1970434; ROM2[9778]<=26'd11123478; ROM3[9778]<=26'd9725621; ROM4[9778]<=26'd23440814;
ROM1[9779]<=26'd1962146; ROM2[9779]<=26'd11112363; ROM3[9779]<=26'd9713976; ROM4[9779]<=26'd23430723;
ROM1[9780]<=26'd1975243; ROM2[9780]<=26'd11117072; ROM3[9780]<=26'd9715799; ROM4[9780]<=26'd23435440;
ROM1[9781]<=26'd1992233; ROM2[9781]<=26'd11125518; ROM3[9781]<=26'd9717878; ROM4[9781]<=26'd23441645;
ROM1[9782]<=26'd1981222; ROM2[9782]<=26'd11113411; ROM3[9782]<=26'd9707406; ROM4[9782]<=26'd23430448;
ROM1[9783]<=26'd1968221; ROM2[9783]<=26'd11106587; ROM3[9783]<=26'd9703500; ROM4[9783]<=26'd23423315;
ROM1[9784]<=26'd1959328; ROM2[9784]<=26'd11105870; ROM3[9784]<=26'd9705660; ROM4[9784]<=26'd23422202;
ROM1[9785]<=26'd1956697; ROM2[9785]<=26'd11106865; ROM3[9785]<=26'd9709725; ROM4[9785]<=26'd23425482;
ROM1[9786]<=26'd1952253; ROM2[9786]<=26'd11108308; ROM3[9786]<=26'd9712284; ROM4[9786]<=26'd23427731;
ROM1[9787]<=26'd1956955; ROM2[9787]<=26'd11112360; ROM3[9787]<=26'd9718064; ROM4[9787]<=26'd23432523;
ROM1[9788]<=26'd1963219; ROM2[9788]<=26'd11110714; ROM3[9788]<=26'd9713753; ROM4[9788]<=26'd23430237;
ROM1[9789]<=26'd1971317; ROM2[9789]<=26'd11110030; ROM3[9789]<=26'd9705907; ROM4[9789]<=26'd23427310;
ROM1[9790]<=26'd1976036; ROM2[9790]<=26'd11111662; ROM3[9790]<=26'd9705450; ROM4[9790]<=26'd23428212;
ROM1[9791]<=26'd1968889; ROM2[9791]<=26'd11109639; ROM3[9791]<=26'd9708157; ROM4[9791]<=26'd23428465;
ROM1[9792]<=26'd1961160; ROM2[9792]<=26'd11110440; ROM3[9792]<=26'd9714133; ROM4[9792]<=26'd23430681;
ROM1[9793]<=26'd1955094; ROM2[9793]<=26'd11108476; ROM3[9793]<=26'd9715928; ROM4[9793]<=26'd23431010;
ROM1[9794]<=26'd1945896; ROM2[9794]<=26'd11104188; ROM3[9794]<=26'd9716614; ROM4[9794]<=26'd23429597;
ROM1[9795]<=26'd1941642; ROM2[9795]<=26'd11102487; ROM3[9795]<=26'd9717748; ROM4[9795]<=26'd23429285;
ROM1[9796]<=26'd1946540; ROM2[9796]<=26'd11102907; ROM3[9796]<=26'd9715833; ROM4[9796]<=26'd23430767;
ROM1[9797]<=26'd1960182; ROM2[9797]<=26'd11105204; ROM3[9797]<=26'd9712358; ROM4[9797]<=26'd23432018;
ROM1[9798]<=26'd1968948; ROM2[9798]<=26'd11103803; ROM3[9798]<=26'd9707781; ROM4[9798]<=26'd23431245;
ROM1[9799]<=26'd1965806; ROM2[9799]<=26'd11101531; ROM3[9799]<=26'd9707568; ROM4[9799]<=26'd23431096;
ROM1[9800]<=26'd1959367; ROM2[9800]<=26'd11100697; ROM3[9800]<=26'd9711916; ROM4[9800]<=26'd23432086;
ROM1[9801]<=26'd1954665; ROM2[9801]<=26'd11101606; ROM3[9801]<=26'd9719348; ROM4[9801]<=26'd23435019;
ROM1[9802]<=26'd1949589; ROM2[9802]<=26'd11101713; ROM3[9802]<=26'd9724773; ROM4[9802]<=26'd23437500;
ROM1[9803]<=26'd1949334; ROM2[9803]<=26'd11104019; ROM3[9803]<=26'd9727771; ROM4[9803]<=26'd23440626;
ROM1[9804]<=26'd1955015; ROM2[9804]<=26'd11106163; ROM3[9804]<=26'd9729235; ROM4[9804]<=26'd23442865;
ROM1[9805]<=26'd1965870; ROM2[9805]<=26'd11106759; ROM3[9805]<=26'd9727522; ROM4[9805]<=26'd23444933;
ROM1[9806]<=26'd1976295; ROM2[9806]<=26'd11104818; ROM3[9806]<=26'd9721396; ROM4[9806]<=26'd23443467;
ROM1[9807]<=26'd1976435; ROM2[9807]<=26'd11104665; ROM3[9807]<=26'd9721228; ROM4[9807]<=26'd23443286;
ROM1[9808]<=26'd1976447; ROM2[9808]<=26'd11109407; ROM3[9808]<=26'd9731649; ROM4[9808]<=26'd23450637;
ROM1[9809]<=26'd1972406; ROM2[9809]<=26'd11111026; ROM3[9809]<=26'd9738269; ROM4[9809]<=26'd23452280;
ROM1[9810]<=26'd1962810; ROM2[9810]<=26'd11105471; ROM3[9810]<=26'd9735484; ROM4[9810]<=26'd23447554;
ROM1[9811]<=26'd1960767; ROM2[9811]<=26'd11107892; ROM3[9811]<=26'd9738327; ROM4[9811]<=26'd23449251;
ROM1[9812]<=26'd1959782; ROM2[9812]<=26'd11109205; ROM3[9812]<=26'd9734462; ROM4[9812]<=26'd23446866;
ROM1[9813]<=26'd1955209; ROM2[9813]<=26'd11099759; ROM3[9813]<=26'd9716924; ROM4[9813]<=26'd23433600;
ROM1[9814]<=26'd1967026; ROM2[9814]<=26'd11103048; ROM3[9814]<=26'd9709923; ROM4[9814]<=26'd23431007;
ROM1[9815]<=26'd1972847; ROM2[9815]<=26'd11107136; ROM3[9815]<=26'd9709872; ROM4[9815]<=26'd23432226;
ROM1[9816]<=26'd1969644; ROM2[9816]<=26'd11110775; ROM3[9816]<=26'd9712872; ROM4[9816]<=26'd23434898;
ROM1[9817]<=26'd1968726; ROM2[9817]<=26'd11116744; ROM3[9817]<=26'd9719804; ROM4[9817]<=26'd23439728;
ROM1[9818]<=26'd1961991; ROM2[9818]<=26'd11115981; ROM3[9818]<=26'd9720648; ROM4[9818]<=26'd23437104;
ROM1[9819]<=26'd1946327; ROM2[9819]<=26'd11105420; ROM3[9819]<=26'd9710488; ROM4[9819]<=26'd23424433;
ROM1[9820]<=26'd1941346; ROM2[9820]<=26'd11099158; ROM3[9820]<=26'd9703784; ROM4[9820]<=26'd23415905;
ROM1[9821]<=26'd1951045; ROM2[9821]<=26'd11103546; ROM3[9821]<=26'd9704825; ROM4[9821]<=26'd23419040;
ROM1[9822]<=26'd1964588; ROM2[9822]<=26'd11107961; ROM3[9822]<=26'd9702535; ROM4[9822]<=26'd23421366;
ROM1[9823]<=26'd1973458; ROM2[9823]<=26'd11111511; ROM3[9823]<=26'd9702012; ROM4[9823]<=26'd23422686;
ROM1[9824]<=26'd1967863; ROM2[9824]<=26'd11110647; ROM3[9824]<=26'd9701721; ROM4[9824]<=26'd23420277;
ROM1[9825]<=26'd1958438; ROM2[9825]<=26'd11109039; ROM3[9825]<=26'd9703666; ROM4[9825]<=26'd23418936;
ROM1[9826]<=26'd1955872; ROM2[9826]<=26'd11110889; ROM3[9826]<=26'd9710005; ROM4[9826]<=26'd23422645;
ROM1[9827]<=26'd1952635; ROM2[9827]<=26'd11111268; ROM3[9827]<=26'd9713817; ROM4[9827]<=26'd23425470;
ROM1[9828]<=26'd1949264; ROM2[9828]<=26'd11109977; ROM3[9828]<=26'd9716901; ROM4[9828]<=26'd23426612;
ROM1[9829]<=26'd1959500; ROM2[9829]<=26'd11115023; ROM3[9829]<=26'd9721672; ROM4[9829]<=26'd23432131;
ROM1[9830]<=26'd1976114; ROM2[9830]<=26'd11121151; ROM3[9830]<=26'd9723019; ROM4[9830]<=26'd23436130;
ROM1[9831]<=26'd1987844; ROM2[9831]<=26'd11121124; ROM3[9831]<=26'd9720232; ROM4[9831]<=26'd23436914;
ROM1[9832]<=26'd1986570; ROM2[9832]<=26'd11118716; ROM3[9832]<=26'd9719842; ROM4[9832]<=26'd23437082;
ROM1[9833]<=26'd1972588; ROM2[9833]<=26'd11110964; ROM3[9833]<=26'd9717477; ROM4[9833]<=26'd23430325;
ROM1[9834]<=26'd1961005; ROM2[9834]<=26'd11106687; ROM3[9834]<=26'd9718125; ROM4[9834]<=26'd23426850;
ROM1[9835]<=26'd1959241; ROM2[9835]<=26'd11108164; ROM3[9835]<=26'd9723541; ROM4[9835]<=26'd23430053;
ROM1[9836]<=26'd1953030; ROM2[9836]<=26'd11106003; ROM3[9836]<=26'd9726586; ROM4[9836]<=26'd23432072;
ROM1[9837]<=26'd1953117; ROM2[9837]<=26'd11105849; ROM3[9837]<=26'd9727780; ROM4[9837]<=26'd23434064;
ROM1[9838]<=26'd1959924; ROM2[9838]<=26'd11105506; ROM3[9838]<=26'd9723543; ROM4[9838]<=26'd23434093;
ROM1[9839]<=26'd1967242; ROM2[9839]<=26'd11100972; ROM3[9839]<=26'd9714231; ROM4[9839]<=26'd23428734;
ROM1[9840]<=26'd1969117; ROM2[9840]<=26'd11096913; ROM3[9840]<=26'd9710330; ROM4[9840]<=26'd23425338;
ROM1[9841]<=26'd1962224; ROM2[9841]<=26'd11095582; ROM3[9841]<=26'd9714328; ROM4[9841]<=26'd23427129;
ROM1[9842]<=26'd1956661; ROM2[9842]<=26'd11096257; ROM3[9842]<=26'd9722555; ROM4[9842]<=26'd23429355;
ROM1[9843]<=26'd1956068; ROM2[9843]<=26'd11098046; ROM3[9843]<=26'd9728412; ROM4[9843]<=26'd23431291;
ROM1[9844]<=26'd1949932; ROM2[9844]<=26'd11097060; ROM3[9844]<=26'd9729855; ROM4[9844]<=26'd23432246;
ROM1[9845]<=26'd1947954; ROM2[9845]<=26'd11097444; ROM3[9845]<=26'd9730288; ROM4[9845]<=26'd23431596;
ROM1[9846]<=26'd1959440; ROM2[9846]<=26'd11103793; ROM3[9846]<=26'd9732756; ROM4[9846]<=26'd23436703;
ROM1[9847]<=26'd1966250; ROM2[9847]<=26'd11102342; ROM3[9847]<=26'd9725939; ROM4[9847]<=26'd23435905;
ROM1[9848]<=26'd1966022; ROM2[9848]<=26'd11095065; ROM3[9848]<=26'd9716609; ROM4[9848]<=26'd23426884;
ROM1[9849]<=26'd1964536; ROM2[9849]<=26'd11093796; ROM3[9849]<=26'd9718417; ROM4[9849]<=26'd23426726;
ROM1[9850]<=26'd1957858; ROM2[9850]<=26'd11092292; ROM3[9850]<=26'd9720971; ROM4[9850]<=26'd23427274;
ROM1[9851]<=26'd1953261; ROM2[9851]<=26'd11093597; ROM3[9851]<=26'd9726519; ROM4[9851]<=26'd23429073;
ROM1[9852]<=26'd1952021; ROM2[9852]<=26'd11098827; ROM3[9852]<=26'd9732596; ROM4[9852]<=26'd23433875;
ROM1[9853]<=26'd1945064; ROM2[9853]<=26'd11097177; ROM3[9853]<=26'd9731077; ROM4[9853]<=26'd23430389;
ROM1[9854]<=26'd1942297; ROM2[9854]<=26'd11093516; ROM3[9854]<=26'd9726732; ROM4[9854]<=26'd23426594;
ROM1[9855]<=26'd1953332; ROM2[9855]<=26'd11094671; ROM3[9855]<=26'd9723865; ROM4[9855]<=26'd23426637;
ROM1[9856]<=26'd1970164; ROM2[9856]<=26'd11100776; ROM3[9856]<=26'd9723510; ROM4[9856]<=26'd23430290;
ROM1[9857]<=26'd1976523; ROM2[9857]<=26'd11106696; ROM3[9857]<=26'd9727112; ROM4[9857]<=26'd23436303;
ROM1[9858]<=26'd1966916; ROM2[9858]<=26'd11102369; ROM3[9858]<=26'd9725075; ROM4[9858]<=26'd23432333;
ROM1[9859]<=26'd1954961; ROM2[9859]<=26'd11096487; ROM3[9859]<=26'd9723040; ROM4[9859]<=26'd23428529;
ROM1[9860]<=26'd1947152; ROM2[9860]<=26'd11093918; ROM3[9860]<=26'd9721074; ROM4[9860]<=26'd23426195;
ROM1[9861]<=26'd1935465; ROM2[9861]<=26'd11088998; ROM3[9861]<=26'd9717894; ROM4[9861]<=26'd23420414;
ROM1[9862]<=26'd1937027; ROM2[9862]<=26'd11090022; ROM3[9862]<=26'd9719819; ROM4[9862]<=26'd23420917;
ROM1[9863]<=26'd1951535; ROM2[9863]<=26'd11097029; ROM3[9863]<=26'd9720388; ROM4[9863]<=26'd23424757;
ROM1[9864]<=26'd1971437; ROM2[9864]<=26'd11104800; ROM3[9864]<=26'd9721805; ROM4[9864]<=26'd23431613;
ROM1[9865]<=26'd1982330; ROM2[9865]<=26'd11109412; ROM3[9865]<=26'd9725946; ROM4[9865]<=26'd23437881;
ROM1[9866]<=26'd1973478; ROM2[9866]<=26'd11104460; ROM3[9866]<=26'd9726214; ROM4[9866]<=26'd23435677;
ROM1[9867]<=26'd1961034; ROM2[9867]<=26'd11099168; ROM3[9867]<=26'd9726544; ROM4[9867]<=26'd23432830;
ROM1[9868]<=26'd1953741; ROM2[9868]<=26'd11096789; ROM3[9868]<=26'd9727518; ROM4[9868]<=26'd23429907;
ROM1[9869]<=26'd1949738; ROM2[9869]<=26'd11096474; ROM3[9869]<=26'd9731903; ROM4[9869]<=26'd23431480;
ROM1[9870]<=26'd1948305; ROM2[9870]<=26'd11096124; ROM3[9870]<=26'd9731994; ROM4[9870]<=26'd23432451;
ROM1[9871]<=26'd1951488; ROM2[9871]<=26'd11093126; ROM3[9871]<=26'd9726247; ROM4[9871]<=26'd23428896;
ROM1[9872]<=26'd1961117; ROM2[9872]<=26'd11090875; ROM3[9872]<=26'd9719379; ROM4[9872]<=26'd23426590;
ROM1[9873]<=26'd1965667; ROM2[9873]<=26'd11090045; ROM3[9873]<=26'd9711990; ROM4[9873]<=26'd23425184;
ROM1[9874]<=26'd1964157; ROM2[9874]<=26'd11093820; ROM3[9874]<=26'd9716118; ROM4[9874]<=26'd23429578;
ROM1[9875]<=26'd1960933; ROM2[9875]<=26'd11097509; ROM3[9875]<=26'd9724355; ROM4[9875]<=26'd23434206;
ROM1[9876]<=26'd1954045; ROM2[9876]<=26'd11096101; ROM3[9876]<=26'd9728038; ROM4[9876]<=26'd23433813;
ROM1[9877]<=26'd1943360; ROM2[9877]<=26'd11091449; ROM3[9877]<=26'd9727626; ROM4[9877]<=26'd23430291;
ROM1[9878]<=26'd1939124; ROM2[9878]<=26'd11091463; ROM3[9878]<=26'd9728034; ROM4[9878]<=26'd23429852;
ROM1[9879]<=26'd1942741; ROM2[9879]<=26'd11093089; ROM3[9879]<=26'd9728744; ROM4[9879]<=26'd23430976;
ROM1[9880]<=26'd1952008; ROM2[9880]<=26'd11094058; ROM3[9880]<=26'd9723778; ROM4[9880]<=26'd23429875;
ROM1[9881]<=26'd1965617; ROM2[9881]<=26'd11097203; ROM3[9881]<=26'd9719006; ROM4[9881]<=26'd23430376;
ROM1[9882]<=26'd1968924; ROM2[9882]<=26'd11101038; ROM3[9882]<=26'd9723276; ROM4[9882]<=26'd23435244;
ROM1[9883]<=26'd1963704; ROM2[9883]<=26'd11102769; ROM3[9883]<=26'd9728796; ROM4[9883]<=26'd23438190;
ROM1[9884]<=26'd1961904; ROM2[9884]<=26'd11108350; ROM3[9884]<=26'd9738223; ROM4[9884]<=26'd23445200;
ROM1[9885]<=26'd1959937; ROM2[9885]<=26'd11112361; ROM3[9885]<=26'd9743289; ROM4[9885]<=26'd23447955;
ROM1[9886]<=26'd1948189; ROM2[9886]<=26'd11105321; ROM3[9886]<=26'd9737087; ROM4[9886]<=26'd23439272;
ROM1[9887]<=26'd1945418; ROM2[9887]<=26'd11103065; ROM3[9887]<=26'd9733746; ROM4[9887]<=26'd23436510;
ROM1[9888]<=26'd1951703; ROM2[9888]<=26'd11104120; ROM3[9888]<=26'd9729553; ROM4[9888]<=26'd23436005;
ROM1[9889]<=26'd1965431; ROM2[9889]<=26'd11104481; ROM3[9889]<=26'd9724617; ROM4[9889]<=26'd23434804;
ROM1[9890]<=26'd1974323; ROM2[9890]<=26'd11108014; ROM3[9890]<=26'd9725276; ROM4[9890]<=26'd23438366;
ROM1[9891]<=26'd1969577; ROM2[9891]<=26'd11111397; ROM3[9891]<=26'd9728325; ROM4[9891]<=26'd23441709;
ROM1[9892]<=26'd1962648; ROM2[9892]<=26'd11112498; ROM3[9892]<=26'd9732534; ROM4[9892]<=26'd23441699;
ROM1[9893]<=26'd1958424; ROM2[9893]<=26'd11111970; ROM3[9893]<=26'd9735123; ROM4[9893]<=26'd23441853;
ROM1[9894]<=26'd1953635; ROM2[9894]<=26'd11111423; ROM3[9894]<=26'd9736869; ROM4[9894]<=26'd23441691;
ROM1[9895]<=26'd1953964; ROM2[9895]<=26'd11114314; ROM3[9895]<=26'd9738882; ROM4[9895]<=26'd23442571;
ROM1[9896]<=26'd1960221; ROM2[9896]<=26'd11115398; ROM3[9896]<=26'd9734037; ROM4[9896]<=26'd23440762;
ROM1[9897]<=26'd1967102; ROM2[9897]<=26'd11112953; ROM3[9897]<=26'd9725947; ROM4[9897]<=26'd23436431;
ROM1[9898]<=26'd1972180; ROM2[9898]<=26'd11112448; ROM3[9898]<=26'd9719180; ROM4[9898]<=26'd23431959;
ROM1[9899]<=26'd1967443; ROM2[9899]<=26'd11109580; ROM3[9899]<=26'd9716772; ROM4[9899]<=26'd23428693;
ROM1[9900]<=26'd1960742; ROM2[9900]<=26'd11107812; ROM3[9900]<=26'd9721039; ROM4[9900]<=26'd23429848;
ROM1[9901]<=26'd1956206; ROM2[9901]<=26'd11109322; ROM3[9901]<=26'd9723449; ROM4[9901]<=26'd23429778;
ROM1[9902]<=26'd1952769; ROM2[9902]<=26'd11112629; ROM3[9902]<=26'd9727997; ROM4[9902]<=26'd23432153;
ROM1[9903]<=26'd1951524; ROM2[9903]<=26'd11114757; ROM3[9903]<=26'd9731971; ROM4[9903]<=26'd23434720;
ROM1[9904]<=26'd1953483; ROM2[9904]<=26'd11114072; ROM3[9904]<=26'd9731590; ROM4[9904]<=26'd23434645;
ROM1[9905]<=26'd1958164; ROM2[9905]<=26'd11109834; ROM3[9905]<=26'd9724912; ROM4[9905]<=26'd23431012;
ROM1[9906]<=26'd1969559; ROM2[9906]<=26'd11109306; ROM3[9906]<=26'd9719548; ROM4[9906]<=26'd23429952;
ROM1[9907]<=26'd1971904; ROM2[9907]<=26'd11110221; ROM3[9907]<=26'd9721402; ROM4[9907]<=26'd23431835;
ROM1[9908]<=26'd1966310; ROM2[9908]<=26'd11108722; ROM3[9908]<=26'd9722865; ROM4[9908]<=26'd23430758;
ROM1[9909]<=26'd1973864; ROM2[9909]<=26'd11120271; ROM3[9909]<=26'd9736667; ROM4[9909]<=26'd23443812;
ROM1[9910]<=26'd1975362; ROM2[9910]<=26'd11124631; ROM3[9910]<=26'd9744735; ROM4[9910]<=26'd23449224;
ROM1[9911]<=26'd1964441; ROM2[9911]<=26'd11118545; ROM3[9911]<=26'd9740243; ROM4[9911]<=26'd23442160;
ROM1[9912]<=26'd1955262; ROM2[9912]<=26'd11111195; ROM3[9912]<=26'd9730166; ROM4[9912]<=26'd23433144;
ROM1[9913]<=26'd1954061; ROM2[9913]<=26'd11103867; ROM3[9913]<=26'd9718701; ROM4[9913]<=26'd23423517;
ROM1[9914]<=26'd1964908; ROM2[9914]<=26'd11104012; ROM3[9914]<=26'd9712828; ROM4[9914]<=26'd23422634;
ROM1[9915]<=26'd1973278; ROM2[9915]<=26'd11107715; ROM3[9915]<=26'd9713558; ROM4[9915]<=26'd23425279;
ROM1[9916]<=26'd1977548; ROM2[9916]<=26'd11116438; ROM3[9916]<=26'd9726031; ROM4[9916]<=26'd23433223;
ROM1[9917]<=26'd1968998; ROM2[9917]<=26'd11115193; ROM3[9917]<=26'd9728914; ROM4[9917]<=26'd23433616;
ROM1[9918]<=26'd1959655; ROM2[9918]<=26'd11110049; ROM3[9918]<=26'd9726115; ROM4[9918]<=26'd23430250;
ROM1[9919]<=26'd1952630; ROM2[9919]<=26'd11107244; ROM3[9919]<=26'd9728064; ROM4[9919]<=26'd23429986;
ROM1[9920]<=26'd1944841; ROM2[9920]<=26'd11101098; ROM3[9920]<=26'd9724544; ROM4[9920]<=26'd23425694;
ROM1[9921]<=26'd1948616; ROM2[9921]<=26'd11100941; ROM3[9921]<=26'd9721599; ROM4[9921]<=26'd23423227;
ROM1[9922]<=26'd1961837; ROM2[9922]<=26'd11104303; ROM3[9922]<=26'd9718813; ROM4[9922]<=26'd23424282;
ROM1[9923]<=26'd1970028; ROM2[9923]<=26'd11106747; ROM3[9923]<=26'd9715171; ROM4[9923]<=26'd23425408;
ROM1[9924]<=26'd1974638; ROM2[9924]<=26'd11113619; ROM3[9924]<=26'd9721872; ROM4[9924]<=26'd23432998;
ROM1[9925]<=26'd1969883; ROM2[9925]<=26'd11112570; ROM3[9925]<=26'd9725555; ROM4[9925]<=26'd23434296;
ROM1[9926]<=26'd1954116; ROM2[9926]<=26'd11102051; ROM3[9926]<=26'd9721512; ROM4[9926]<=26'd23425076;
ROM1[9927]<=26'd1948588; ROM2[9927]<=26'd11099126; ROM3[9927]<=26'd9723414; ROM4[9927]<=26'd23424296;
ROM1[9928]<=26'd1945459; ROM2[9928]<=26'd11099831; ROM3[9928]<=26'd9723998; ROM4[9928]<=26'd23424477;
ROM1[9929]<=26'd1948974; ROM2[9929]<=26'd11104103; ROM3[9929]<=26'd9725785; ROM4[9929]<=26'd23426130;
ROM1[9930]<=26'd1967757; ROM2[9930]<=26'd11114670; ROM3[9930]<=26'd9730589; ROM4[9930]<=26'd23435078;
ROM1[9931]<=26'd1981018; ROM2[9931]<=26'd11117439; ROM3[9931]<=26'd9726653; ROM4[9931]<=26'd23436888;
ROM1[9932]<=26'd1976588; ROM2[9932]<=26'd11111899; ROM3[9932]<=26'd9723574; ROM4[9932]<=26'd23433270;
ROM1[9933]<=26'd1967387; ROM2[9933]<=26'd11107518; ROM3[9933]<=26'd9723503; ROM4[9933]<=26'd23431302;
ROM1[9934]<=26'd1958486; ROM2[9934]<=26'd11104893; ROM3[9934]<=26'd9724255; ROM4[9934]<=26'd23429827;
ROM1[9935]<=26'd1953534; ROM2[9935]<=26'd11104336; ROM3[9935]<=26'd9728688; ROM4[9935]<=26'd23430067;
ROM1[9936]<=26'd1950220; ROM2[9936]<=26'd11106577; ROM3[9936]<=26'd9732172; ROM4[9936]<=26'd23431341;
ROM1[9937]<=26'd1953658; ROM2[9937]<=26'd11108495; ROM3[9937]<=26'd9734188; ROM4[9937]<=26'd23433241;
ROM1[9938]<=26'd1963964; ROM2[9938]<=26'd11110436; ROM3[9938]<=26'd9732220; ROM4[9938]<=26'd23435094;
ROM1[9939]<=26'd1974917; ROM2[9939]<=26'd11111414; ROM3[9939]<=26'd9726542; ROM4[9939]<=26'd23433888;
ROM1[9940]<=26'd1977395; ROM2[9940]<=26'd11109548; ROM3[9940]<=26'd9723839; ROM4[9940]<=26'd23431630;
ROM1[9941]<=26'd1976308; ROM2[9941]<=26'd11114038; ROM3[9941]<=26'd9730705; ROM4[9941]<=26'd23436149;
ROM1[9942]<=26'd1978151; ROM2[9942]<=26'd11122423; ROM3[9942]<=26'd9741044; ROM4[9942]<=26'd23444379;
ROM1[9943]<=26'd1968354; ROM2[9943]<=26'd11116360; ROM3[9943]<=26'd9736482; ROM4[9943]<=26'd23439882;
ROM1[9944]<=26'd1955691; ROM2[9944]<=26'd11110030; ROM3[9944]<=26'd9730870; ROM4[9944]<=26'd23434922;
ROM1[9945]<=26'd1955649; ROM2[9945]<=26'd11112779; ROM3[9945]<=26'd9731760; ROM4[9945]<=26'd23436261;
ROM1[9946]<=26'd1958028; ROM2[9946]<=26'd11111909; ROM3[9946]<=26'd9726888; ROM4[9946]<=26'd23432407;
ROM1[9947]<=26'd1973902; ROM2[9947]<=26'd11119363; ROM3[9947]<=26'd9726233; ROM4[9947]<=26'd23436308;
ROM1[9948]<=26'd1986193; ROM2[9948]<=26'd11122314; ROM3[9948]<=26'd9724793; ROM4[9948]<=26'd23437874;
ROM1[9949]<=26'd1980431; ROM2[9949]<=26'd11117019; ROM3[9949]<=26'd9719751; ROM4[9949]<=26'd23434052;
ROM1[9950]<=26'd1971716; ROM2[9950]<=26'd11116328; ROM3[9950]<=26'd9722289; ROM4[9950]<=26'd23435381;
ROM1[9951]<=26'd1969618; ROM2[9951]<=26'd11119210; ROM3[9951]<=26'd9730213; ROM4[9951]<=26'd23438816;
ROM1[9952]<=26'd1965673; ROM2[9952]<=26'd11117975; ROM3[9952]<=26'd9732882; ROM4[9952]<=26'd23438316;
ROM1[9953]<=26'd1955461; ROM2[9953]<=26'd11111676; ROM3[9953]<=26'd9731308; ROM4[9953]<=26'd23435210;
ROM1[9954]<=26'd1956377; ROM2[9954]<=26'd11109797; ROM3[9954]<=26'd9731482; ROM4[9954]<=26'd23434210;
ROM1[9955]<=26'd1970831; ROM2[9955]<=26'd11113638; ROM3[9955]<=26'd9732687; ROM4[9955]<=26'd23438079;
ROM1[9956]<=26'd1990156; ROM2[9956]<=26'd11123263; ROM3[9956]<=26'd9737816; ROM4[9956]<=26'd23448831;
ROM1[9957]<=26'd1999048; ROM2[9957]<=26'd11132854; ROM3[9957]<=26'd9747988; ROM4[9957]<=26'd23458242;
ROM1[9958]<=26'd1988281; ROM2[9958]<=26'd11127603; ROM3[9958]<=26'd9745315; ROM4[9958]<=26'd23453627;
ROM1[9959]<=26'd1968004; ROM2[9959]<=26'd11114684; ROM3[9959]<=26'd9736758; ROM4[9959]<=26'd23443078;
ROM1[9960]<=26'd1961394; ROM2[9960]<=26'd11112343; ROM3[9960]<=26'd9739933; ROM4[9960]<=26'd23445143;
ROM1[9961]<=26'd1955743; ROM2[9961]<=26'd11109059; ROM3[9961]<=26'd9742485; ROM4[9961]<=26'd23443929;
ROM1[9962]<=26'd1960324; ROM2[9962]<=26'd11112782; ROM3[9962]<=26'd9746752; ROM4[9962]<=26'd23446313;
ROM1[9963]<=26'd1973604; ROM2[9963]<=26'd11118258; ROM3[9963]<=26'd9748156; ROM4[9963]<=26'd23450621;
ROM1[9964]<=26'd1974542; ROM2[9964]<=26'd11107106; ROM3[9964]<=26'd9729973; ROM4[9964]<=26'd23438465;
ROM1[9965]<=26'd1971171; ROM2[9965]<=26'd11099546; ROM3[9965]<=26'd9720400; ROM4[9965]<=26'd23431560;
ROM1[9966]<=26'd1967402; ROM2[9966]<=26'd11099849; ROM3[9966]<=26'd9725443; ROM4[9966]<=26'd23433107;
ROM1[9967]<=26'd1963661; ROM2[9967]<=26'd11103003; ROM3[9967]<=26'd9731001; ROM4[9967]<=26'd23436362;
ROM1[9968]<=26'd1965533; ROM2[9968]<=26'd11108943; ROM3[9968]<=26'd9739667; ROM4[9968]<=26'd23441096;
ROM1[9969]<=26'd1962856; ROM2[9969]<=26'd11110127; ROM3[9969]<=26'd9742183; ROM4[9969]<=26'd23441525;
ROM1[9970]<=26'd1956311; ROM2[9970]<=26'd11107475; ROM3[9970]<=26'd9737143; ROM4[9970]<=26'd23437915;
ROM1[9971]<=26'd1962211; ROM2[9971]<=26'd11107072; ROM3[9971]<=26'd9732995; ROM4[9971]<=26'd23437351;
ROM1[9972]<=26'd1973673; ROM2[9972]<=26'd11108672; ROM3[9972]<=26'd9726445; ROM4[9972]<=26'd23436494;
ROM1[9973]<=26'd1983123; ROM2[9973]<=26'd11113093; ROM3[9973]<=26'd9726099; ROM4[9973]<=26'd23439362;
ROM1[9974]<=26'd1984217; ROM2[9974]<=26'd11115244; ROM3[9974]<=26'd9729534; ROM4[9974]<=26'd23443347;
ROM1[9975]<=26'd1973903; ROM2[9975]<=26'd11113728; ROM3[9975]<=26'd9732680; ROM4[9975]<=26'd23441080;
ROM1[9976]<=26'd1965617; ROM2[9976]<=26'd11113046; ROM3[9976]<=26'd9736502; ROM4[9976]<=26'd23440661;
ROM1[9977]<=26'd1956099; ROM2[9977]<=26'd11109629; ROM3[9977]<=26'd9733662; ROM4[9977]<=26'd23437727;
ROM1[9978]<=26'd1950249; ROM2[9978]<=26'd11108367; ROM3[9978]<=26'd9731812; ROM4[9978]<=26'd23434977;
ROM1[9979]<=26'd1957261; ROM2[9979]<=26'd11112688; ROM3[9979]<=26'd9733748; ROM4[9979]<=26'd23438415;
ROM1[9980]<=26'd1968230; ROM2[9980]<=26'd11115955; ROM3[9980]<=26'd9730204; ROM4[9980]<=26'd23438623;
ROM1[9981]<=26'd1972036; ROM2[9981]<=26'd11109287; ROM3[9981]<=26'd9716701; ROM4[9981]<=26'd23430163;
ROM1[9982]<=26'd1969754; ROM2[9982]<=26'd11106972; ROM3[9982]<=26'd9714074; ROM4[9982]<=26'd23428338;
ROM1[9983]<=26'd1962081; ROM2[9983]<=26'd11105459; ROM3[9983]<=26'd9713752; ROM4[9983]<=26'd23425083;
ROM1[9984]<=26'd1954731; ROM2[9984]<=26'd11101934; ROM3[9984]<=26'd9714814; ROM4[9984]<=26'd23422571;
ROM1[9985]<=26'd1955288; ROM2[9985]<=26'd11106524; ROM3[9985]<=26'd9720818; ROM4[9985]<=26'd23427124;
ROM1[9986]<=26'd1955353; ROM2[9986]<=26'd11110415; ROM3[9986]<=26'd9726347; ROM4[9986]<=26'd23431502;
ROM1[9987]<=26'd1959782; ROM2[9987]<=26'd11112988; ROM3[9987]<=26'd9729007; ROM4[9987]<=26'd23434712;
ROM1[9988]<=26'd1962600; ROM2[9988]<=26'd11108563; ROM3[9988]<=26'd9719690; ROM4[9988]<=26'd23428694;
ROM1[9989]<=26'd1977704; ROM2[9989]<=26'd11111766; ROM3[9989]<=26'd9716670; ROM4[9989]<=26'd23430876;
ROM1[9990]<=26'd1984288; ROM2[9990]<=26'd11111861; ROM3[9990]<=26'd9715474; ROM4[9990]<=26'd23431544;
ROM1[9991]<=26'd1972566; ROM2[9991]<=26'd11106108; ROM3[9991]<=26'd9711152; ROM4[9991]<=26'd23427717;
ROM1[9992]<=26'd1967761; ROM2[9992]<=26'd11109034; ROM3[9992]<=26'd9717622; ROM4[9992]<=26'd23431728;
ROM1[9993]<=26'd1966344; ROM2[9993]<=26'd11111708; ROM3[9993]<=26'd9725679; ROM4[9993]<=26'd23435261;
ROM1[9994]<=26'd1959101; ROM2[9994]<=26'd11110029; ROM3[9994]<=26'd9726985; ROM4[9994]<=26'd23434599;
ROM1[9995]<=26'd1956274; ROM2[9995]<=26'd11107493; ROM3[9995]<=26'd9726255; ROM4[9995]<=26'd23432165;
ROM1[9996]<=26'd1964079; ROM2[9996]<=26'd11110395; ROM3[9996]<=26'd9726822; ROM4[9996]<=26'd23435261;
ROM1[9997]<=26'd1977698; ROM2[9997]<=26'd11115119; ROM3[9997]<=26'd9725560; ROM4[9997]<=26'd23438485;
ROM1[9998]<=26'd1988271; ROM2[9998]<=26'd11117073; ROM3[9998]<=26'd9724014; ROM4[9998]<=26'd23440717;
ROM1[9999]<=26'd1985939; ROM2[9999]<=26'd11116688; ROM3[9999]<=26'd9726915; ROM4[9999]<=26'd23441133;


	end
	else begin
		if(cnt == 127) begin
				cnt<=0;
			end
		//원래는 addr이다.
		data1 <= ROM1[cnt];
		data2 <= ROM2[cnt];
		data3 <= ROM3[cnt];
		data4 <= ROM4[cnt];
		cnt <= cnt+1;
	end
end
endmodule 
