/*
 * MUL2
 * have to consider input sequence
 */

module ONE_UNIT_MUL3 (
    input clk_mul,
    input en_mul,

    // z
    input signed [25:0] zi1, zi2, zi3, zi4,
    // zTw
    input signed [25:0] zw1_11, zw1_12, zw1_13, zw1_14,
    input signed [25:0] zw1_21, zw1_22, zw1_23, zw1_24,
    input signed [25:0] zw1_31, zw1_32, zw1_33, zw1_34,
    input signed [25:0] zw1_41, zw1_42, zw1_43, zw1_44,

    input signed [25:0] zw2_11, zw2_12, zw2_13, zw2_14,
    input signed [25:0] zw2_21, zw2_22, zw2_23, zw2_24,
    input signed [25:0] zw2_31, zw2_32, zw2_33, zw2_34,
    input signed [25:0] zw2_41, zw2_42, zw2_43, zw2_44,

    input signed [25:0] zw3_11, zw3_12, zw3_13, zw3_14,
    input signed [25:0] zw3_21, zw3_22, zw3_23, zw3_24,
    input signed [25:0] zw3_31, zw3_32, zw3_33, zw3_34,
    input signed [25:0] zw3_41, zw3_42, zw3_43, zw3_44,

    input signed [25:0] zw4_11, zw4_12, zw4_13, zw4_14,
    input signed [25:0] zw4_21, zw4_22, zw4_23, zw4_24,
    input signed [25:0] zw4_31, zw4_32, zw4_33, zw4_34,
    input signed [25:0] zw4_41, zw4_42, zw4_43, zw4_44,
    // (zTw)^2
    input signed [25:0] i1_11, i1_12, i1_13, i1_14,
    input signed [25:0] i1_21, i1_22, i1_23, i1_24,
    input signed [25:0] i1_31, i1_32, i1_33, i1_34,
    input signed [25:0] i1_41, i1_42, i1_43, i1_44,

    input signed [25:0] i2_11, i2_12, i2_13, i2_14,
    input signed [25:0] i2_21, i2_22, i2_23, i2_24,
    input signed [25:0] i2_31, i2_32, i2_33, i2_34,
    input signed [25:0] i2_41, i2_42, i2_43, i2_44,

    input signed [25:0] i3_11, i3_12, i3_13, i3_14,
    input signed [25:0] i3_21, i3_22, i3_23, i3_24,
    input signed [25:0] i3_31, i3_32, i3_33, i3_34,
    input signed [25:0] i3_41, i3_42, i3_43, i3_44,

    input signed [25:0] i4_11, i4_12, i4_13, i4_14,
    input signed [25:0] i4_21, i4_22, i4_23, i4_24,
    input signed [25:0] i4_31, i4_32, i4_33, i4_34,
    input signed [25:0] i4_41, i4_42, i4_43, i4_44,
    
    // z
    output reg signed [25:0] zo1, zo2, zo3, zo4,

    // (zTw)^2
    output signed [25:0] zTw_3_1_11, zTw_3_1_12, zTw_3_1_13, zTw_3_1_14,
    output signed [25:0] zTw_3_1_21, zTw_3_1_22, zTw_3_1_23, zTw_3_1_24,
    output signed [25:0] zTw_3_1_31, zTw_3_1_32, zTw_3_1_33, zTw_3_1_34,
    output signed [25:0] zTw_3_1_41, zTw_3_1_42, zTw_3_1_43, zTw_3_1_44,

    output signed [25:0] zTw_3_2_11, zTw_3_2_12, zTw_3_2_13, zTw_3_2_14,
    output signed [25:0] zTw_3_2_21, zTw_3_2_22, zTw_3_2_23, zTw_3_2_24,
    output signed [25:0] zTw_3_2_31, zTw_3_2_32, zTw_3_2_33, zTw_3_2_34,
    output signed [25:0] zTw_3_2_41, zTw_3_2_42, zTw_3_2_43, zTw_3_2_44,

    output signed [25:0] zTw_3_3_11, zTw_3_3_12, zTw_3_3_13, zTw_3_3_14,
    output signed [25:0] zTw_3_3_21, zTw_3_3_22, zTw_3_3_23, zTw_3_3_24,
    output signed [25:0] zTw_3_3_31, zTw_3_3_32, zTw_3_3_33, zTw_3_3_34,
    output signed [25:0] zTw_3_3_41, zTw_3_3_42, zTw_3_3_43, zTw_3_3_44,

    output signed [25:0] zTw_3_4_11, zTw_3_4_12, zTw_3_4_13, zTw_3_4_14,
    output signed [25:0] zTw_3_4_21, zTw_3_4_22, zTw_3_4_23, zTw_3_4_24,
    output signed [25:0] zTw_3_4_31, zTw_3_4_32, zTw_3_4_33, zTw_3_4_34,
    output signed [25:0] zTw_3_4_41, zTw_3_4_42, zTw_3_4_43, zTw_3_4_44
);

reg signed [51:0] zTw_3_1_11_reg, zTw_3_1_12_reg, zTw_3_1_13_reg, zTw_3_1_14_reg;
reg signed [51:0] zTw_3_1_21_reg, zTw_3_1_22_reg, zTw_3_1_23_reg, zTw_3_1_24_reg;
reg signed [51:0] zTw_3_1_31_reg, zTw_3_1_32_reg, zTw_3_1_33_reg, zTw_3_1_34_reg;
reg signed [51:0] zTw_3_1_41_reg, zTw_3_1_42_reg, zTw_3_1_43_reg, zTw_3_1_44_reg;

reg signed [51:0] zTw_3_2_11_reg, zTw_3_2_12_reg, zTw_3_2_13_reg, zTw_3_2_14_reg;
reg signed [51:0] zTw_3_2_21_reg, zTw_3_2_22_reg, zTw_3_2_23_reg, zTw_3_2_24_reg;
reg signed [51:0] zTw_3_2_31_reg, zTw_3_2_32_reg, zTw_3_2_33_reg, zTw_3_2_34_reg;
reg signed [51:0] zTw_3_2_41_reg, zTw_3_2_42_reg, zTw_3_2_43_reg, zTw_3_2_44_reg;

reg signed [51:0] zTw_3_3_11_reg, zTw_3_3_12_reg, zTw_3_3_13_reg, zTw_3_3_14_reg;
reg signed [51:0] zTw_3_3_21_reg, zTw_3_3_22_reg, zTw_3_3_23_reg, zTw_3_3_24_reg;
reg signed [51:0] zTw_3_3_31_reg, zTw_3_3_32_reg, zTw_3_3_33_reg, zTw_3_3_34_reg;
reg signed [51:0] zTw_3_3_41_reg, zTw_3_3_42_reg, zTw_3_3_43_reg, zTw_3_3_44_reg;

reg signed [51:0] zTw_3_4_11_reg, zTw_3_4_12_reg, zTw_3_4_13_reg, zTw_3_4_14_reg;
reg signed [51:0] zTw_3_4_21_reg, zTw_3_4_22_reg, zTw_3_4_23_reg, zTw_3_4_24_reg;
reg signed [51:0] zTw_3_4_31_reg, zTw_3_4_32_reg, zTw_3_4_33_reg, zTw_3_4_34_reg;
reg signed [51:0] zTw_3_4_41_reg, zTw_3_4_42_reg, zTw_3_4_43_reg, zTw_3_4_44_reg;

assign zTw_3_1_11 = zTw_3_1_11_reg[38:13];
assign zTw_3_1_12 = zTw_3_1_12_reg[38:13];
assign zTw_3_1_13 = zTw_3_1_13_reg[38:13];
assign zTw_3_1_14 = zTw_3_1_14_reg[38:13];
assign zTw_3_1_21 = zTw_3_1_21_reg[38:13];
assign zTw_3_1_22 = zTw_3_1_22_reg[38:13];
assign zTw_3_1_23 = zTw_3_1_23_reg[38:13];
assign zTw_3_1_24 = zTw_3_1_24_reg[38:13];
assign zTw_3_1_31 = zTw_3_1_31_reg[38:13];
assign zTw_3_1_32 = zTw_3_1_32_reg[38:13];
assign zTw_3_1_33 = zTw_3_1_33_reg[38:13];
assign zTw_3_1_34 = zTw_3_1_34_reg[38:13];
assign zTw_3_1_41 = zTw_3_1_41_reg[38:13];
assign zTw_3_1_42 = zTw_3_1_42_reg[38:13];
assign zTw_3_1_43 = zTw_3_1_43_reg[38:13];
assign zTw_3_1_44 = zTw_3_1_44_reg[38:13];

assign zTw_3_2_11 = zTw_3_2_11_reg[38:13];
assign zTw_3_2_12 = zTw_3_2_12_reg[38:13];
assign zTw_3_2_13 = zTw_3_2_13_reg[38:13];
assign zTw_3_2_14 = zTw_3_2_14_reg[38:13];
assign zTw_3_2_21 = zTw_3_2_21_reg[38:13];
assign zTw_3_2_22 = zTw_3_2_22_reg[38:13];
assign zTw_3_2_23 = zTw_3_2_23_reg[38:13];
assign zTw_3_2_24 = zTw_3_2_24_reg[38:13];
assign zTw_3_2_31 = zTw_3_2_31_reg[38:13];
assign zTw_3_2_32 = zTw_3_2_32_reg[38:13];
assign zTw_3_2_33 = zTw_3_2_33_reg[38:13];
assign zTw_3_2_34 = zTw_3_2_34_reg[38:13];
assign zTw_3_2_41 = zTw_3_2_41_reg[38:13];
assign zTw_3_2_42 = zTw_3_2_42_reg[38:13];
assign zTw_3_2_43 = zTw_3_2_43_reg[38:13];
assign zTw_3_2_44 = zTw_3_2_44_reg[38:13];

assign zTw_3_3_11 = zTw_3_3_11_reg[38:13];
assign zTw_3_3_12 = zTw_3_3_12_reg[38:13];
assign zTw_3_3_13 = zTw_3_3_13_reg[38:13];
assign zTw_3_3_14 = zTw_3_3_14_reg[38:13];
assign zTw_3_3_21 = zTw_3_3_21_reg[38:13];
assign zTw_3_3_22 = zTw_3_3_22_reg[38:13];
assign zTw_3_3_23 = zTw_3_3_23_reg[38:13];
assign zTw_3_3_24 = zTw_3_3_24_reg[38:13];
assign zTw_3_3_31 = zTw_3_3_31_reg[38:13];
assign zTw_3_3_32 = zTw_3_3_32_reg[38:13];
assign zTw_3_3_33 = zTw_3_3_33_reg[38:13];
assign zTw_3_3_34 = zTw_3_3_34_reg[38:13];
assign zTw_3_3_41 = zTw_3_3_41_reg[38:13];
assign zTw_3_3_42 = zTw_3_3_42_reg[38:13];
assign zTw_3_3_43 = zTw_3_3_43_reg[38:13];
assign zTw_3_3_44 = zTw_3_3_44_reg[38:13];

assign zTw_3_4_11 = zTw_3_4_11_reg[38:13];
assign zTw_3_4_12 = zTw_3_4_12_reg[38:13];
assign zTw_3_4_13 = zTw_3_4_13_reg[38:13];
assign zTw_3_4_14 = zTw_3_4_14_reg[38:13];
assign zTw_3_4_21 = zTw_3_4_21_reg[38:13];
assign zTw_3_4_22 = zTw_3_4_22_reg[38:13];
assign zTw_3_4_23 = zTw_3_4_23_reg[38:13];
assign zTw_3_4_24 = zTw_3_4_24_reg[38:13];
assign zTw_3_4_31 = zTw_3_4_31_reg[38:13];
assign zTw_3_4_32 = zTw_3_4_32_reg[38:13];
assign zTw_3_4_33 = zTw_3_4_33_reg[38:13];
assign zTw_3_4_34 = zTw_3_4_34_reg[38:13];
assign zTw_3_4_41 = zTw_3_4_41_reg[38:13];
assign zTw_3_4_42 = zTw_3_4_42_reg[38:13];
assign zTw_3_4_43 = zTw_3_4_43_reg[38:13];
assign zTw_3_4_44 = zTw_3_4_44_reg[38:13];

always @(posedge clk_mul)
begin
    zo1 <= zi1;
    zo2 <= zi2;
    zo3 <= zi3;
    zo4 <= zi4;
    if (en_mul) begin
        // active
        zTw_3_1_11_reg <= zw1_11 * i1_11 + zw1_12 * i1_21 + zw1_13 * i1_31 + zw1_14 * i1_41;
        zTw_3_1_12_reg <= zw1_11 * i1_12 + zw1_12 * i1_22 + zw1_13 * i1_32 + zw1_14 * i1_42;
        zTw_3_1_13_reg <= zw1_11 * i1_13 + zw1_12 * i1_23 + zw1_13 * i1_33 + zw1_14 * i1_43;
        zTw_3_1_14_reg <= zw1_11 * i1_14 + zw1_12 * i1_24 + zw1_13 * i1_34 + zw1_14 * i1_44;
        zTw_3_1_21_reg <= zw1_21 * i1_11 + zw1_22 * i1_21 + zw1_23 * i1_31 + zw1_24 * i1_41;
        zTw_3_1_22_reg <= zw1_21 * i1_12 + zw1_22 * i1_22 + zw1_23 * i1_32 + zw1_24 * i1_42;
        zTw_3_1_23_reg <= zw1_21 * i1_13 + zw1_22 * i1_23 + zw1_23 * i1_33 + zw1_24 * i1_43;
        zTw_3_1_24_reg <= zw1_21 * i1_14 + zw1_22 * i1_24 + zw1_23 * i1_34 + zw1_24 * i1_44;
        zTw_3_1_31_reg <= zw1_31 * i1_11 + zw1_32 * i1_21 + zw1_33 * i1_31 + zw1_34 * i1_41;
        zTw_3_1_32_reg <= zw1_31 * i1_12 + zw1_32 * i1_22 + zw1_33 * i1_32 + zw1_34 * i1_42;
        zTw_3_1_33_reg <= zw1_31 * i1_13 + zw1_32 * i1_23 + zw1_33 * i1_33 + zw1_34 * i1_43;
        zTw_3_1_34_reg <= zw1_31 * i1_14 + zw1_32 * i1_24 + zw1_33 * i1_34 + zw1_34 * i1_44;
        zTw_3_1_41_reg <= zw1_41 * i1_11 + zw1_42 * i1_21 + zw1_43 * i1_31 + zw1_44 * i1_41;
        zTw_3_1_42_reg <= zw1_41 * i1_12 + zw1_42 * i1_22 + zw1_43 * i1_32 + zw1_44 * i1_42;
        zTw_3_1_43_reg <= zw1_41 * i1_13 + zw1_42 * i1_23 + zw1_43 * i1_33 + zw1_44 * i1_43;
        zTw_3_1_44_reg <= zw1_41 * i1_14 + zw1_42 * i1_24 + zw1_43 * i1_34 + zw1_44 * i1_44;

        zTw_3_2_11_reg <= zw2_11 * i2_11 + zw2_12 * i2_21 + zw2_13 * i2_31 + zw2_14 * i2_41;
        zTw_3_2_12_reg <= zw2_11 * i2_12 + zw2_12 * i2_22 + zw2_13 * i2_32 + zw2_14 * i2_42;
        zTw_3_2_13_reg <= zw2_11 * i2_13 + zw2_12 * i2_23 + zw2_13 * i2_33 + zw2_14 * i2_43;
        zTw_3_2_14_reg <= zw2_11 * i2_14 + zw2_12 * i2_24 + zw2_13 * i2_34 + zw2_14 * i2_44;
        zTw_3_2_21_reg <= zw2_21 * i2_11 + zw2_22 * i2_21 + zw2_23 * i2_31 + zw2_24 * i2_41;
        zTw_3_2_22_reg <= zw2_21 * i2_12 + zw2_22 * i2_22 + zw2_23 * i2_32 + zw2_24 * i2_42;
        zTw_3_2_23_reg <= zw2_21 * i2_13 + zw2_22 * i2_23 + zw2_23 * i2_33 + zw2_24 * i2_43;
        zTw_3_2_24_reg <= zw2_21 * i2_14 + zw2_22 * i2_24 + zw2_23 * i2_34 + zw2_24 * i2_44;
        zTw_3_2_31_reg <= zw2_31 * i2_11 + zw2_32 * i2_21 + zw2_33 * i2_31 + zw2_34 * i2_41;
        zTw_3_2_32_reg <= zw2_31 * i2_12 + zw2_32 * i2_22 + zw2_33 * i2_32 + zw2_34 * i2_42;
        zTw_3_2_33_reg <= zw2_31 * i2_13 + zw2_32 * i2_23 + zw2_33 * i2_33 + zw2_34 * i2_43;
        zTw_3_2_34_reg <= zw2_31 * i2_14 + zw2_32 * i2_24 + zw2_33 * i2_34 + zw2_34 * i2_44;
        zTw_3_2_41_reg <= zw2_41 * i2_11 + zw2_42 * i2_21 + zw2_43 * i2_31 + zw2_44 * i2_41;
        zTw_3_2_42_reg <= zw2_41 * i2_12 + zw2_42 * i2_22 + zw2_43 * i2_32 + zw2_44 * i2_42;
        zTw_3_2_43_reg <= zw2_41 * i2_13 + zw2_42 * i2_23 + zw2_43 * i2_33 + zw2_44 * i2_43;
        zTw_3_2_44_reg <= zw2_41 * i2_14 + zw2_42 * i2_24 + zw2_43 * i2_34 + zw2_44 * i2_44;

        zTw_3_3_11_reg <= zw3_11 * i3_11 + zw3_12 * i3_21 + zw3_13 * i3_31 + zw3_14 * i3_41;
        zTw_3_3_12_reg <= zw3_11 * i3_12 + zw3_12 * i3_22 + zw3_13 * i3_32 + zw3_14 * i3_42;
        zTw_3_3_13_reg <= zw3_11 * i3_13 + zw3_12 * i3_23 + zw3_13 * i3_33 + zw3_14 * i3_43;
        zTw_3_3_14_reg <= zw3_11 * i3_14 + zw3_12 * i3_24 + zw3_13 * i3_34 + zw3_14 * i3_44;
        zTw_3_3_21_reg <= zw3_21 * i3_11 + zw3_22 * i3_21 + zw3_23 * i3_31 + zw3_24 * i3_41;
        zTw_3_3_22_reg <= zw3_21 * i3_12 + zw3_22 * i3_22 + zw3_23 * i3_32 + zw3_24 * i3_42;
        zTw_3_3_23_reg <= zw3_21 * i3_13 + zw3_22 * i3_23 + zw3_23 * i3_33 + zw3_24 * i3_43;
        zTw_3_3_24_reg <= zw3_21 * i3_14 + zw3_22 * i3_24 + zw3_23 * i3_34 + zw3_24 * i3_44;
        zTw_3_3_31_reg <= zw3_31 * i3_11 + zw3_32 * i3_21 + zw3_33 * i3_31 + zw3_34 * i3_41;
        zTw_3_3_32_reg <= zw3_31 * i3_12 + zw3_32 * i3_22 + zw3_33 * i3_32 + zw3_34 * i3_42;
        zTw_3_3_33_reg <= zw3_31 * i3_13 + zw3_32 * i3_23 + zw3_33 * i3_33 + zw3_34 * i3_43;
        zTw_3_3_34_reg <= zw3_31 * i3_14 + zw3_32 * i3_24 + zw3_33 * i3_34 + zw3_34 * i3_44;
        zTw_3_3_41_reg <= zw3_41 * i3_11 + zw3_42 * i3_21 + zw3_43 * i3_31 + zw3_44 * i3_41;
        zTw_3_3_42_reg <= zw3_41 * i3_12 + zw3_42 * i3_22 + zw3_43 * i3_32 + zw3_44 * i3_42;
        zTw_3_3_43_reg <= zw3_41 * i3_13 + zw3_42 * i3_23 + zw3_43 * i3_33 + zw3_44 * i3_43;
        zTw_3_3_44_reg <= zw3_41 * i3_14 + zw3_42 * i3_24 + zw3_43 * i3_34 + zw3_44 * i3_44;

        zTw_3_4_11_reg <= zw4_11 * i4_11 + zw4_12 * i4_21 + zw4_13 * i4_31 + zw4_14 * i4_41;
        zTw_3_4_12_reg <= zw4_11 * i4_12 + zw4_12 * i4_22 + zw4_13 * i4_32 + zw4_14 * i4_42;
        zTw_3_4_13_reg <= zw4_11 * i4_13 + zw4_12 * i4_23 + zw4_13 * i4_33 + zw4_14 * i4_43;
        zTw_3_4_14_reg <= zw4_11 * i4_14 + zw4_12 * i4_24 + zw4_13 * i4_34 + zw4_14 * i4_44;
        zTw_3_4_21_reg <= zw4_21 * i4_11 + zw4_22 * i4_21 + zw4_23 * i4_31 + zw4_24 * i4_41;
        zTw_3_4_22_reg <= zw4_21 * i4_12 + zw4_22 * i4_22 + zw4_23 * i4_32 + zw4_24 * i4_42;
        zTw_3_4_23_reg <= zw4_21 * i4_13 + zw4_22 * i4_23 + zw4_23 * i4_33 + zw4_24 * i4_43;
        zTw_3_4_24_reg <= zw4_21 * i4_14 + zw4_22 * i4_24 + zw4_23 * i4_34 + zw4_24 * i4_44;
        zTw_3_4_31_reg <= zw4_31 * i4_11 + zw4_32 * i4_21 + zw4_33 * i4_31 + zw4_34 * i4_41;
        zTw_3_4_32_reg <= zw4_31 * i4_12 + zw4_32 * i4_22 + zw4_33 * i4_32 + zw4_34 * i4_42;
        zTw_3_4_33_reg <= zw4_31 * i4_13 + zw4_32 * i4_23 + zw4_33 * i4_33 + zw4_34 * i4_43;
        zTw_3_4_34_reg <= zw4_31 * i4_14 + zw4_32 * i4_24 + zw4_33 * i4_34 + zw4_34 * i4_44;
        zTw_3_4_41_reg <= zw4_41 * i4_11 + zw4_42 * i4_21 + zw4_43 * i4_31 + zw4_44 * i4_41;
        zTw_3_4_42_reg <= zw4_41 * i4_12 + zw4_42 * i4_22 + zw4_43 * i4_32 + zw4_44 * i4_42;
        zTw_3_4_43_reg <= zw4_41 * i4_13 + zw4_42 * i4_23 + zw4_43 * i4_33 + zw4_44 * i4_43;
        zTw_3_4_44_reg <= zw4_41 * i4_14 + zw4_42 * i4_24 + zw4_43 * i4_34 + zw4_44 * i4_44;
    end else begin
        // zTw_3_1_11_reg <= i1_11;
        // zTw_3_1_12_reg <= i1_12;
        // zTw_3_1_13_reg <= i1_13;
        // zTw_3_1_14_reg <= i1_14;
        // zTw_3_1_21_reg <= i1_21;
        // zTw_3_1_22_reg <= i1_22;
        // zTw_3_1_23_reg <= i1_23;
        // zTw_3_1_24_reg <= i1_24;
        // zTw_3_1_31_reg <= i1_31;
        // zTw_3_1_32_reg <= i1_32;
        // zTw_3_1_33_reg <= i1_33;
        // zTw_3_1_34_reg <= i1_34;
        // zTw_3_1_41_reg <= i1_41;
        // zTw_3_1_42_reg <= i1_42;
        // zTw_3_1_43_reg <= i1_43;
        // zTw_3_1_44_reg <= i1_44;

        // zTw_3_2_11_reg <= i2_11;
        // zTw_3_2_12_reg <= i2_12;
        // zTw_3_2_13_reg <= i2_13;
        // zTw_3_2_14_reg <= i2_14;
        // zTw_3_2_21_reg <= i2_21;
        // zTw_3_2_22_reg <= i2_22;
        // zTw_3_2_23_reg <= i2_23;
        // zTw_3_2_24_reg <= i2_24;
        // zTw_3_2_31_reg <= i2_31;
        // zTw_3_2_32_reg <= i2_32;
        // zTw_3_2_33_reg <= i2_33;
        // zTw_3_2_34_reg <= i2_34;
        // zTw_3_2_41_reg <= i2_41;
        // zTw_3_2_42_reg <= i2_42;
        // zTw_3_2_43_reg <= i2_43;
        // zTw_3_2_44_reg <= i2_44;

        // zTw_3_3_11_reg <= i3_11;
        // zTw_3_3_12_reg <= i3_12;
        // zTw_3_3_13_reg <= i3_13;
        // zTw_3_3_14_reg <= i3_14;
        // zTw_3_3_21_reg <= i3_21;
        // zTw_3_3_22_reg <= i3_22;
        // zTw_3_3_23_reg <= i3_23;
        // zTw_3_3_24_reg <= i3_24;
        // zTw_3_3_31_reg <= i3_31;
        // zTw_3_3_32_reg <= i3_32;
        // zTw_3_3_33_reg <= i3_33;
        // zTw_3_3_34_reg <= i3_34;
        // zTw_3_3_41_reg <= i3_41;
        // zTw_3_3_42_reg <= i3_42;
        // zTw_3_3_43_reg <= i3_43;
        // zTw_3_3_44_reg <= i3_44;

        // zTw_3_4_11_reg <= i4_11;
        // zTw_3_4_12_reg <= i4_12;
        // zTw_3_4_13_reg <= i4_13;
        // zTw_3_4_14_reg <= i4_14;
        // zTw_3_4_21_reg <= i4_21;
        // zTw_3_4_22_reg <= i4_22;
        // zTw_3_4_23_reg <= i4_23;
        // zTw_3_4_24_reg <= i4_24;
        // zTw_3_4_31_reg <= i4_31;
        // zTw_3_4_32_reg <= i4_32;
        // zTw_3_4_33_reg <= i4_33;
        // zTw_3_4_34_reg <= i4_34;
        // zTw_3_4_41_reg <= i4_41;
        // zTw_3_4_42_reg <= i4_42;
        // zTw_3_4_43_reg <= i4_43;
        // zTw_3_4_44_reg <= i4_44;
    end
end
    
endmodule