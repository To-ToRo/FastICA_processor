module Multiplier(
X11,X12,X13,X14,
X21,X22,X23,X24,
X31,X32,X33,X34,
X41,X42,X43,X44,
Y11,Y12,Y13,Y14,
Y21,Y22,Y23,Y24,
Y31,Y32,Y33,Y34,
Y41,Y42,Y43,Y44,
Z11,Z12,Z13,Z14,
Z21,Z22,Z23,Z24,
Z31,Z32,Z33,Z34,
Z41,Z42,Z43,Z44);

input signed [63:0] X11,X12,X13,X14,X21,X22,X23,X24,X31,X32,X33,X34,X41,X42,X43,X44;
input signed [63:0] Y11,Y12,Y13,Y14,Y21,Y22,Y23,Y24,Y31,Y32,Y33,Y34,Y41,Y42,Y43,Y44;
output wire signed [63:0] Z11,Z12,Z13,Z14,Z21,Z22,Z23,Z24,Z31,Z32,Z33,Z34,Z41,Z42,Z43,Z44;

wire signed [127:0] XY11,XY12,XY13,XY14,XY21,XY22,XY23,XY24,XY31,XY32,XY33,XY34,XY41,XY42,XY43,XY44;

assign XY11 = X11*Y11 + X12*Y21 + X13*Y31 + X14*Y41;
assign XY12 = X11*Y12 + X12*Y22 + X13*Y32 + X14*Y42;
assign XY13 = X11*Y13 + X12*Y23 + X13*Y33 + X14*Y43;
assign XY14 = X11*Y14 + X12*Y24 + X13*Y34 + X14*Y44;
assign XY21 = X21*Y11 + X22*Y21 + X23*Y31 + X24*Y41;
assign XY22 = X21*Y12 + X22*Y22 + X23*Y32 + X24*Y42;
assign XY23 = X21*Y13 + X22*Y23 + X23*Y33 + X24*Y43;
assign XY24 = X21*Y14 + X22*Y24 + X23*Y34 + X24*Y44;
assign XY31 = X31*Y11 + X32*Y21 + X33*Y31 + X34*Y41;
assign XY32 = X31*Y12 + X32*Y22 + X33*Y32 + X34*Y42;
assign XY33 = X31*Y13 + X32*Y23 + X33*Y33 + X34*Y43;
assign XY34 = X31*Y14 + X32*Y24 + X33*Y34 + X34*Y44;
assign XY41 = X41*Y11 + X42*Y21 + X43*Y31 + X44*Y41;
assign XY42 = X41*Y12 + X42*Y22 + X43*Y32 + X44*Y42;
assign XY43 = X41*Y13 + X42*Y23 + X43*Y33 + X44*Y43;
assign XY44 = X41*Y14 + X42*Y24 + X43*Y34 + X44*Y44;

assign Z11 = XY11[95:32];
assign Z12 = XY12[95:32];
assign Z13 = XY13[95:32];
assign Z14 = XY14[95:32];
assign Z21 = XY21[95:32];
assign Z22 = XY22[95:32];
assign Z23 = XY23[95:32];
assign Z24 = XY24[95:32];
assign Z31 = XY31[95:32];
assign Z32 = XY32[95:32];
assign Z33 = XY33[95:32];
assign Z34 = XY34[95:32];
assign Z41 = XY41[95:32];
assign Z42 = XY42[95:32];
assign Z43 = XY43[95:32];
assign Z44 = XY44[95:32];

endmodule