//출처 : https://verilogguide.readthedocs.io/en/latest/verilog/designs.html#read-only-memory-rom

module ROM(
    input wire clk,
	input wire En,
    input wire  [13:0] addr,
    output reg signed [15:0] data1,
	output reg signed [15:0] data2,
	output reg signed [15:0] data3,
	output reg signed [15:0] data4
);

//ROM[0]의 크기 : 16bit(한 시그널의 크기) * 4(4개의 시그널) 
// 각각의 시그널이 총 1000sample이 있으므로 addr은  16비트로 표현(0~39999 < 0~65536) 

reg unsigned [16:0] ROM1[0:9999];
reg unsigned [16:0] ROM2[0:9999];
reg unsigned [16:0] ROM3[0:9999];
reg unsigned [16:0] ROM4[0:9999];
reg [6:0] cnt;

always @(posedge clk) begin
	if(!En) begin
		cnt<=0;
ROM1[0]<=16'd4788; ROM2[0]<=16'd0; ROM3[0]<=16'd23830; ROM4[0]<=16'd57282;
ROM1[1]<=16'd4790; ROM2[1]<=16'd0; ROM3[1]<=16'd23840; ROM4[1]<=16'd57289;
ROM1[2]<=16'd4765; ROM2[2]<=16'd0; ROM3[2]<=16'd23839; ROM4[2]<=16'd57287;
ROM1[3]<=16'd4730; ROM2[3]<=16'd0; ROM3[3]<=16'd23824; ROM4[3]<=16'd57266;
ROM1[4]<=16'd4717; ROM2[4]<=16'd0; ROM3[4]<=16'd23823; ROM4[4]<=16'd57264;
ROM1[5]<=16'd4706; ROM2[5]<=16'd0; ROM3[5]<=16'd23827; ROM4[5]<=16'd57263;
ROM1[6]<=16'd4717; ROM2[6]<=16'd0; ROM3[6]<=16'd23837; ROM4[6]<=16'd57272;
ROM1[7]<=16'd4734; ROM2[7]<=16'd0; ROM3[7]<=16'd23821; ROM4[7]<=16'd57267;
ROM1[8]<=16'd4743; ROM2[8]<=16'd0; ROM3[8]<=16'd23789; ROM4[8]<=16'd57247;
ROM1[9]<=16'd4756; ROM2[9]<=16'd0; ROM3[9]<=16'd23787; ROM4[9]<=16'd57251;
ROM1[10]<=16'd4744; ROM2[10]<=16'd0; ROM3[10]<=16'd23794; ROM4[10]<=16'd57254;
ROM1[11]<=16'd4736; ROM2[11]<=16'd0; ROM3[11]<=16'd23813; ROM4[11]<=16'd57265;
ROM1[12]<=16'd4727; ROM2[12]<=16'd0; ROM3[12]<=16'd23823; ROM4[12]<=16'd57271;
ROM1[13]<=16'd4700; ROM2[13]<=16'd0; ROM3[13]<=16'd23818; ROM4[13]<=16'd57263;
ROM1[14]<=16'd4687; ROM2[14]<=16'd0; ROM3[14]<=16'd23813; ROM4[14]<=16'd57251;
ROM1[15]<=16'd4706; ROM2[15]<=16'd0; ROM3[15]<=16'd23807; ROM4[15]<=16'd57252;
ROM1[16]<=16'd4756; ROM2[16]<=16'd0; ROM3[16]<=16'd23814; ROM4[16]<=16'd57270;
ROM1[17]<=16'd4785; ROM2[17]<=16'd0; ROM3[17]<=16'd23814; ROM4[17]<=16'd57281;
ROM1[18]<=16'd4762; ROM2[18]<=16'd0; ROM3[18]<=16'd23792; ROM4[18]<=16'd57263;
ROM1[19]<=16'd4730; ROM2[19]<=16'd0; ROM3[19]<=16'd23787; ROM4[19]<=16'd57251;
ROM1[20]<=16'd4713; ROM2[20]<=16'd0; ROM3[20]<=16'd23792; ROM4[20]<=16'd57244;
ROM1[21]<=16'd4696; ROM2[21]<=16'd0; ROM3[21]<=16'd23786; ROM4[21]<=16'd57230;
ROM1[22]<=16'd4685; ROM2[22]<=16'd0; ROM3[22]<=16'd23791; ROM4[22]<=16'd57236;
ROM1[23]<=16'd4695; ROM2[23]<=16'd0; ROM3[23]<=16'd23790; ROM4[23]<=16'd57241;
ROM1[24]<=16'd4718; ROM2[24]<=16'd0; ROM3[24]<=16'd23774; ROM4[24]<=16'd57233;
ROM1[25]<=16'd4745; ROM2[25]<=16'd0; ROM3[25]<=16'd23757; ROM4[25]<=16'd57232;
ROM1[26]<=16'd4748; ROM2[26]<=16'd0; ROM3[26]<=16'd23758; ROM4[26]<=16'd57235;
ROM1[27]<=16'd4733; ROM2[27]<=16'd0; ROM3[27]<=16'd23764; ROM4[27]<=16'd57234;
ROM1[28]<=16'd4711; ROM2[28]<=16'd0; ROM3[28]<=16'd23772; ROM4[28]<=16'd57233;
ROM1[29]<=16'd4691; ROM2[29]<=16'd0; ROM3[29]<=16'd23774; ROM4[29]<=16'd57230;
ROM1[30]<=16'd4680; ROM2[30]<=16'd0; ROM3[30]<=16'd23774; ROM4[30]<=16'd57230;
ROM1[31]<=16'd4692; ROM2[31]<=16'd0; ROM3[31]<=16'd23779; ROM4[31]<=16'd57235;
ROM1[32]<=16'd4724; ROM2[32]<=16'd0; ROM3[32]<=16'd23777; ROM4[32]<=16'd57244;
ROM1[33]<=16'd4759; ROM2[33]<=16'd0; ROM3[33]<=16'd23770; ROM4[33]<=16'd57252;
ROM1[34]<=16'd4765; ROM2[34]<=16'd0; ROM3[34]<=16'd23776; ROM4[34]<=16'd57258;
ROM1[35]<=16'd4750; ROM2[35]<=16'd0; ROM3[35]<=16'd23789; ROM4[35]<=16'd57265;
ROM1[36]<=16'd4739; ROM2[36]<=16'd0; ROM3[36]<=16'd23805; ROM4[36]<=16'd57271;
ROM1[37]<=16'd4735; ROM2[37]<=16'd0; ROM3[37]<=16'd23818; ROM4[37]<=16'd57270;
ROM1[38]<=16'd4733; ROM2[38]<=16'd0; ROM3[38]<=16'd23827; ROM4[38]<=16'd57272;
ROM1[39]<=16'd4728; ROM2[39]<=16'd0; ROM3[39]<=16'd23826; ROM4[39]<=16'd57268;
ROM1[40]<=16'd4744; ROM2[40]<=16'd0; ROM3[40]<=16'd23825; ROM4[40]<=16'd57271;
ROM1[41]<=16'd4759; ROM2[41]<=16'd0; ROM3[41]<=16'd23799; ROM4[41]<=16'd57257;
ROM1[42]<=16'd4763; ROM2[42]<=16'd0; ROM3[42]<=16'd23775; ROM4[42]<=16'd57242;
ROM1[43]<=16'd4757; ROM2[43]<=16'd0; ROM3[43]<=16'd23779; ROM4[43]<=16'd57241;
ROM1[44]<=16'd4740; ROM2[44]<=16'd0; ROM3[44]<=16'd23786; ROM4[44]<=16'd57240;
ROM1[45]<=16'd4720; ROM2[45]<=16'd0; ROM3[45]<=16'd23792; ROM4[45]<=16'd57244;
ROM1[46]<=16'd4709; ROM2[46]<=16'd0; ROM3[46]<=16'd23796; ROM4[46]<=16'd57243;
ROM1[47]<=16'd4701; ROM2[47]<=16'd0; ROM3[47]<=16'd23795; ROM4[47]<=16'd57240;
ROM1[48]<=16'd4711; ROM2[48]<=16'd0; ROM3[48]<=16'd23797; ROM4[48]<=16'd57246;
ROM1[49]<=16'd4738; ROM2[49]<=16'd0; ROM3[49]<=16'd23790; ROM4[49]<=16'd57249;
ROM1[50]<=16'd4758; ROM2[50]<=16'd0; ROM3[50]<=16'd23778; ROM4[50]<=16'd57242;
ROM1[51]<=16'd4766; ROM2[51]<=16'd0; ROM3[51]<=16'd23789; ROM4[51]<=16'd57256;
ROM1[52]<=16'd4743; ROM2[52]<=16'd0; ROM3[52]<=16'd23786; ROM4[52]<=16'd57254;
ROM1[53]<=16'd4713; ROM2[53]<=16'd0; ROM3[53]<=16'd23775; ROM4[53]<=16'd57233;
ROM1[54]<=16'd4710; ROM2[54]<=16'd0; ROM3[54]<=16'd23788; ROM4[54]<=16'd57239;
ROM1[55]<=16'd4700; ROM2[55]<=16'd0; ROM3[55]<=16'd23798; ROM4[55]<=16'd57243;
ROM1[56]<=16'd4695; ROM2[56]<=16'd0; ROM3[56]<=16'd23792; ROM4[56]<=16'd57235;
ROM1[57]<=16'd4723; ROM2[57]<=16'd0; ROM3[57]<=16'd23791; ROM4[57]<=16'd57240;
ROM1[58]<=16'd4758; ROM2[58]<=16'd0; ROM3[58]<=16'd23781; ROM4[58]<=16'd57242;
ROM1[59]<=16'd4762; ROM2[59]<=16'd0; ROM3[59]<=16'd23772; ROM4[59]<=16'd57241;
ROM1[60]<=16'd4749; ROM2[60]<=16'd0; ROM3[60]<=16'd23781; ROM4[60]<=16'd57244;
ROM1[61]<=16'd4748; ROM2[61]<=16'd0; ROM3[61]<=16'd23811; ROM4[61]<=16'd57266;
ROM1[62]<=16'd4752; ROM2[62]<=16'd0; ROM3[62]<=16'd23838; ROM4[62]<=16'd57288;
ROM1[63]<=16'd4728; ROM2[63]<=16'd0; ROM3[63]<=16'd23834; ROM4[63]<=16'd57274;
ROM1[64]<=16'd4714; ROM2[64]<=16'd0; ROM3[64]<=16'd23826; ROM4[64]<=16'd57265;
ROM1[65]<=16'd4728; ROM2[65]<=16'd0; ROM3[65]<=16'd23822; ROM4[65]<=16'd57265;
ROM1[66]<=16'd4752; ROM2[66]<=16'd0; ROM3[66]<=16'd23806; ROM4[66]<=16'd57261;
ROM1[67]<=16'd4772; ROM2[67]<=16'd0; ROM3[67]<=16'd23800; ROM4[67]<=16'd57266;
ROM1[68]<=16'd4770; ROM2[68]<=16'd0; ROM3[68]<=16'd23807; ROM4[68]<=16'd57270;
ROM1[69]<=16'd4751; ROM2[69]<=16'd0; ROM3[69]<=16'd23815; ROM4[69]<=16'd57269;
ROM1[70]<=16'd4734; ROM2[70]<=16'd0; ROM3[70]<=16'd23824; ROM4[70]<=16'd57269;
ROM1[71]<=16'd4733; ROM2[71]<=16'd0; ROM3[71]<=16'd23840; ROM4[71]<=16'd57279;
ROM1[72]<=16'd4730; ROM2[72]<=16'd0; ROM3[72]<=16'd23848; ROM4[72]<=16'd57284;
ROM1[73]<=16'd4734; ROM2[73]<=16'd0; ROM3[73]<=16'd23838; ROM4[73]<=16'd57281;
ROM1[74]<=16'd4748; ROM2[74]<=16'd0; ROM3[74]<=16'd23813; ROM4[74]<=16'd57269;
ROM1[75]<=16'd4760; ROM2[75]<=16'd0; ROM3[75]<=16'd23782; ROM4[75]<=16'd57249;
ROM1[76]<=16'd4751; ROM2[76]<=16'd0; ROM3[76]<=16'd23769; ROM4[76]<=16'd57237;
ROM1[77]<=16'd4739; ROM2[77]<=16'd0; ROM3[77]<=16'd23780; ROM4[77]<=16'd57245;
ROM1[78]<=16'd4735; ROM2[78]<=16'd0; ROM3[78]<=16'd23803; ROM4[78]<=16'd57262;
ROM1[79]<=16'd4712; ROM2[79]<=16'd0; ROM3[79]<=16'd23801; ROM4[79]<=16'd57252;
ROM1[80]<=16'd4695; ROM2[80]<=16'd0; ROM3[80]<=16'd23798; ROM4[80]<=16'd57248;
ROM1[81]<=16'd4691; ROM2[81]<=16'd0; ROM3[81]<=16'd23791; ROM4[81]<=16'd57245;
ROM1[82]<=16'd4702; ROM2[82]<=16'd0; ROM3[82]<=16'd23766; ROM4[82]<=16'd57225;
ROM1[83]<=16'd4733; ROM2[83]<=16'd0; ROM3[83]<=16'd23752; ROM4[83]<=16'd57224;
ROM1[84]<=16'd4744; ROM2[84]<=16'd0; ROM3[84]<=16'd23755; ROM4[84]<=16'd57232;
ROM1[85]<=16'd4736; ROM2[85]<=16'd0; ROM3[85]<=16'd23765; ROM4[85]<=16'd57237;
ROM1[86]<=16'd4717; ROM2[86]<=16'd0; ROM3[86]<=16'd23769; ROM4[86]<=16'd57233;
ROM1[87]<=16'd4711; ROM2[87]<=16'd0; ROM3[87]<=16'd23777; ROM4[87]<=16'd57237;
ROM1[88]<=16'd4698; ROM2[88]<=16'd0; ROM3[88]<=16'd23787; ROM4[88]<=16'd57239;
ROM1[89]<=16'd4680; ROM2[89]<=16'd0; ROM3[89]<=16'd23775; ROM4[89]<=16'd57222;
ROM1[90]<=16'd4694; ROM2[90]<=16'd0; ROM3[90]<=16'd23773; ROM4[90]<=16'd57225;
ROM1[91]<=16'd4727; ROM2[91]<=16'd0; ROM3[91]<=16'd23766; ROM4[91]<=16'd57233;
ROM1[92]<=16'd4735; ROM2[92]<=16'd0; ROM3[92]<=16'd23746; ROM4[92]<=16'd57219;
ROM1[93]<=16'd4729; ROM2[93]<=16'd0; ROM3[93]<=16'd23747; ROM4[93]<=16'd57220;
ROM1[94]<=16'd4718; ROM2[94]<=16'd0; ROM3[94]<=16'd23764; ROM4[94]<=16'd57230;
ROM1[95]<=16'd4689; ROM2[95]<=16'd0; ROM3[95]<=16'd23759; ROM4[95]<=16'd57219;
ROM1[96]<=16'd4680; ROM2[96]<=16'd0; ROM3[96]<=16'd23770; ROM4[96]<=16'd57225;
ROM1[97]<=16'd4689; ROM2[97]<=16'd0; ROM3[97]<=16'd23795; ROM4[97]<=16'd57243;
ROM1[98]<=16'd4702; ROM2[98]<=16'd0; ROM3[98]<=16'd23795; ROM4[98]<=16'd57248;
ROM1[99]<=16'd4716; ROM2[99]<=16'd0; ROM3[99]<=16'd23777; ROM4[99]<=16'd57239;
ROM1[100]<=16'd4731; ROM2[100]<=16'd0; ROM3[100]<=16'd23752; ROM4[100]<=16'd57225;
ROM1[101]<=16'd4721; ROM2[101]<=16'd0; ROM3[101]<=16'd23742; ROM4[101]<=16'd57217;
ROM1[102]<=16'd4696; ROM2[102]<=16'd0; ROM3[102]<=16'd23737; ROM4[102]<=16'd57208;
ROM1[103]<=16'd4691; ROM2[103]<=16'd0; ROM3[103]<=16'd23755; ROM4[103]<=16'd57214;
ROM1[104]<=16'd4692; ROM2[104]<=16'd0; ROM3[104]<=16'd23767; ROM4[104]<=16'd57224;
ROM1[105]<=16'd4676; ROM2[105]<=16'd0; ROM3[105]<=16'd23765; ROM4[105]<=16'd57218;
ROM1[106]<=16'd4682; ROM2[106]<=16'd0; ROM3[106]<=16'd23764; ROM4[106]<=16'd57215;
ROM1[107]<=16'd4715; ROM2[107]<=16'd0; ROM3[107]<=16'd23769; ROM4[107]<=16'd57231;
ROM1[108]<=16'd4753; ROM2[108]<=16'd0; ROM3[108]<=16'd23770; ROM4[108]<=16'd57243;
ROM1[109]<=16'd4758; ROM2[109]<=16'd0; ROM3[109]<=16'd23766; ROM4[109]<=16'd57244;
ROM1[110]<=16'd4746; ROM2[110]<=16'd0; ROM3[110]<=16'd23773; ROM4[110]<=16'd57248;
ROM1[111]<=16'd4734; ROM2[111]<=16'd0; ROM3[111]<=16'd23786; ROM4[111]<=16'd57251;
ROM1[112]<=16'd4731; ROM2[112]<=16'd0; ROM3[112]<=16'd23806; ROM4[112]<=16'd57261;
ROM1[113]<=16'd4719; ROM2[113]<=16'd0; ROM3[113]<=16'd23813; ROM4[113]<=16'd57263;
ROM1[114]<=16'd4702; ROM2[114]<=16'd0; ROM3[114]<=16'd23802; ROM4[114]<=16'd57252;
ROM1[115]<=16'd4710; ROM2[115]<=16'd0; ROM3[115]<=16'd23793; ROM4[115]<=16'd57245;
ROM1[116]<=16'd4741; ROM2[116]<=16'd0; ROM3[116]<=16'd23782; ROM4[116]<=16'd57240;
ROM1[117]<=16'd4772; ROM2[117]<=16'd0; ROM3[117]<=16'd23780; ROM4[117]<=16'd57245;
ROM1[118]<=16'd4780; ROM2[118]<=16'd0; ROM3[118]<=16'd23797; ROM4[118]<=16'd57260;
ROM1[119]<=16'd4763; ROM2[119]<=16'd0; ROM3[119]<=16'd23807; ROM4[119]<=16'd57267;
ROM1[120]<=16'd4744; ROM2[120]<=16'd0; ROM3[120]<=16'd23811; ROM4[120]<=16'd57271;
ROM1[121]<=16'd4734; ROM2[121]<=16'd0; ROM3[121]<=16'd23824; ROM4[121]<=16'd57278;
ROM1[122]<=16'd4748; ROM2[122]<=16'd0; ROM3[122]<=16'd23848; ROM4[122]<=16'd57298;
ROM1[123]<=16'd4759; ROM2[123]<=16'd0; ROM3[123]<=16'd23838; ROM4[123]<=16'd57298;
ROM1[124]<=16'd4764; ROM2[124]<=16'd0; ROM3[124]<=16'd23799; ROM4[124]<=16'd57269;
ROM1[125]<=16'd4775; ROM2[125]<=16'd0; ROM3[125]<=16'd23769; ROM4[125]<=16'd57254;
ROM1[126]<=16'd4760; ROM2[126]<=16'd0; ROM3[126]<=16'd23759; ROM4[126]<=16'd57247;
ROM1[127]<=16'd4752; ROM2[127]<=16'd0; ROM3[127]<=16'd23776; ROM4[127]<=16'd57252;
ROM1[128]<=16'd4738; ROM2[128]<=16'd0; ROM3[128]<=16'd23791; ROM4[128]<=16'd57259;
ROM1[129]<=16'd4721; ROM2[129]<=16'd0; ROM3[129]<=16'd23795; ROM4[129]<=16'd57256;
ROM1[130]<=16'd4703; ROM2[130]<=16'd0; ROM3[130]<=16'd23795; ROM4[130]<=16'd57247;
ROM1[131]<=16'd4700; ROM2[131]<=16'd0; ROM3[131]<=16'd23795; ROM4[131]<=16'd57244;
ROM1[132]<=16'd4724; ROM2[132]<=16'd0; ROM3[132]<=16'd23795; ROM4[132]<=16'd57248;
ROM1[133]<=16'd4754; ROM2[133]<=16'd0; ROM3[133]<=16'd23790; ROM4[133]<=16'd57255;
ROM1[134]<=16'd4764; ROM2[134]<=16'd0; ROM3[134]<=16'd23789; ROM4[134]<=16'd57258;
ROM1[135]<=16'd4747; ROM2[135]<=16'd0; ROM3[135]<=16'd23794; ROM4[135]<=16'd57256;
ROM1[136]<=16'd4719; ROM2[136]<=16'd0; ROM3[136]<=16'd23793; ROM4[136]<=16'd57246;
ROM1[137]<=16'd4699; ROM2[137]<=16'd0; ROM3[137]<=16'd23790; ROM4[137]<=16'd57234;
ROM1[138]<=16'd4666; ROM2[138]<=16'd0; ROM3[138]<=16'd23784; ROM4[138]<=16'd57222;
ROM1[139]<=16'd4657; ROM2[139]<=16'd0; ROM3[139]<=16'd23781; ROM4[139]<=16'd57219;
ROM1[140]<=16'd4688; ROM2[140]<=16'd0; ROM3[140]<=16'd23789; ROM4[140]<=16'd57237;
ROM1[141]<=16'd4749; ROM2[141]<=16'd0; ROM3[141]<=16'd23805; ROM4[141]<=16'd57269;
ROM1[142]<=16'd4777; ROM2[142]<=16'd0; ROM3[142]<=16'd23806; ROM4[142]<=16'd57281;
ROM1[143]<=16'd4752; ROM2[143]<=16'd0; ROM3[143]<=16'd23791; ROM4[143]<=16'd57263;
ROM1[144]<=16'd4725; ROM2[144]<=16'd0; ROM3[144]<=16'd23786; ROM4[144]<=16'd57254;
ROM1[145]<=16'd4686; ROM2[145]<=16'd0; ROM3[145]<=16'd23770; ROM4[145]<=16'd57228;
ROM1[146]<=16'd4658; ROM2[146]<=16'd0; ROM3[146]<=16'd23760; ROM4[146]<=16'd57210;
ROM1[147]<=16'd4654; ROM2[147]<=16'd0; ROM3[147]<=16'd23765; ROM4[147]<=16'd57214;
ROM1[148]<=16'd4659; ROM2[148]<=16'd0; ROM3[148]<=16'd23762; ROM4[148]<=16'd57215;
ROM1[149]<=16'd4683; ROM2[149]<=16'd0; ROM3[149]<=16'd23747; ROM4[149]<=16'd57213;
ROM1[150]<=16'd4706; ROM2[150]<=16'd0; ROM3[150]<=16'd23729; ROM4[150]<=16'd57202;
ROM1[151]<=16'd4707; ROM2[151]<=16'd0; ROM3[151]<=16'd23737; ROM4[151]<=16'd57206;
ROM1[152]<=16'd4692; ROM2[152]<=16'd0; ROM3[152]<=16'd23750; ROM4[152]<=16'd57209;
ROM1[153]<=16'd4666; ROM2[153]<=16'd0; ROM3[153]<=16'd23754; ROM4[153]<=16'd57203;
ROM1[154]<=16'd4658; ROM2[154]<=16'd0; ROM3[154]<=16'd23766; ROM4[154]<=16'd57214;
ROM1[155]<=16'd4658; ROM2[155]<=16'd0; ROM3[155]<=16'd23783; ROM4[155]<=16'd57221;
ROM1[156]<=16'd4671; ROM2[156]<=16'd0; ROM3[156]<=16'd23789; ROM4[156]<=16'd57227;
ROM1[157]<=16'd4709; ROM2[157]<=16'd0; ROM3[157]<=16'd23793; ROM4[157]<=16'd57240;
ROM1[158]<=16'd4741; ROM2[158]<=16'd0; ROM3[158]<=16'd23780; ROM4[158]<=16'd57233;
ROM1[159]<=16'd4742; ROM2[159]<=16'd0; ROM3[159]<=16'd23766; ROM4[159]<=16'd57227;
ROM1[160]<=16'd4727; ROM2[160]<=16'd0; ROM3[160]<=16'd23768; ROM4[160]<=16'd57226;
ROM1[161]<=16'd4707; ROM2[161]<=16'd0; ROM3[161]<=16'd23772; ROM4[161]<=16'd57225;
ROM1[162]<=16'd4694; ROM2[162]<=16'd0; ROM3[162]<=16'd23775; ROM4[162]<=16'd57227;
ROM1[163]<=16'd4689; ROM2[163]<=16'd0; ROM3[163]<=16'd23789; ROM4[163]<=16'd57232;
ROM1[164]<=16'd4691; ROM2[164]<=16'd0; ROM3[164]<=16'd23795; ROM4[164]<=16'd57237;
ROM1[165]<=16'd4712; ROM2[165]<=16'd0; ROM3[165]<=16'd23790; ROM4[165]<=16'd57238;
ROM1[166]<=16'd4743; ROM2[166]<=16'd0; ROM3[166]<=16'd23785; ROM4[166]<=16'd57238;
ROM1[167]<=16'd4755; ROM2[167]<=16'd0; ROM3[167]<=16'd23768; ROM4[167]<=16'd57232;
ROM1[168]<=16'd4753; ROM2[168]<=16'd0; ROM3[168]<=16'd23777; ROM4[168]<=16'd57239;
ROM1[169]<=16'd4740; ROM2[169]<=16'd0; ROM3[169]<=16'd23787; ROM4[169]<=16'd57240;
ROM1[170]<=16'd4712; ROM2[170]<=16'd0; ROM3[170]<=16'd23777; ROM4[170]<=16'd57226;
ROM1[171]<=16'd4693; ROM2[171]<=16'd0; ROM3[171]<=16'd23773; ROM4[171]<=16'd57221;
ROM1[172]<=16'd4686; ROM2[172]<=16'd0; ROM3[172]<=16'd23776; ROM4[172]<=16'd57219;
ROM1[173]<=16'd4709; ROM2[173]<=16'd0; ROM3[173]<=16'd23786; ROM4[173]<=16'd57235;
ROM1[174]<=16'd4747; ROM2[174]<=16'd0; ROM3[174]<=16'd23783; ROM4[174]<=16'd57238;
ROM1[175]<=16'd4771; ROM2[175]<=16'd0; ROM3[175]<=16'd23769; ROM4[175]<=16'd57234;
ROM1[176]<=16'd4763; ROM2[176]<=16'd0; ROM3[176]<=16'd23759; ROM4[176]<=16'd57230;
ROM1[177]<=16'd4736; ROM2[177]<=16'd0; ROM3[177]<=16'd23758; ROM4[177]<=16'd57223;
ROM1[178]<=16'd4721; ROM2[178]<=16'd0; ROM3[178]<=16'd23771; ROM4[178]<=16'd57231;
ROM1[179]<=16'd4712; ROM2[179]<=16'd0; ROM3[179]<=16'd23783; ROM4[179]<=16'd57241;
ROM1[180]<=16'd4700; ROM2[180]<=16'd0; ROM3[180]<=16'd23790; ROM4[180]<=16'd57240;
ROM1[181]<=16'd4700; ROM2[181]<=16'd0; ROM3[181]<=16'd23783; ROM4[181]<=16'd57229;
ROM1[182]<=16'd4729; ROM2[182]<=16'd0; ROM3[182]<=16'd23778; ROM4[182]<=16'd57237;
ROM1[183]<=16'd4773; ROM2[183]<=16'd0; ROM3[183]<=16'd23779; ROM4[183]<=16'd57249;
ROM1[184]<=16'd4776; ROM2[184]<=16'd0; ROM3[184]<=16'd23774; ROM4[184]<=16'd57248;
ROM1[185]<=16'd4746; ROM2[185]<=16'd0; ROM3[185]<=16'd23765; ROM4[185]<=16'd57241;
ROM1[186]<=16'd4720; ROM2[186]<=16'd0; ROM3[186]<=16'd23771; ROM4[186]<=16'd57239;
ROM1[187]<=16'd4703; ROM2[187]<=16'd0; ROM3[187]<=16'd23776; ROM4[187]<=16'd57238;
ROM1[188]<=16'd4706; ROM2[188]<=16'd0; ROM3[188]<=16'd23796; ROM4[188]<=16'd57253;
ROM1[189]<=16'd4711; ROM2[189]<=16'd0; ROM3[189]<=16'd23813; ROM4[189]<=16'd57261;
ROM1[190]<=16'd4701; ROM2[190]<=16'd0; ROM3[190]<=16'd23789; ROM4[190]<=16'd57242;
ROM1[191]<=16'd4724; ROM2[191]<=16'd0; ROM3[191]<=16'd23771; ROM4[191]<=16'd57235;
ROM1[192]<=16'd4742; ROM2[192]<=16'd0; ROM3[192]<=16'd23761; ROM4[192]<=16'd57233;
ROM1[193]<=16'd4729; ROM2[193]<=16'd0; ROM3[193]<=16'd23756; ROM4[193]<=16'd57231;
ROM1[194]<=16'd4727; ROM2[194]<=16'd0; ROM3[194]<=16'd23778; ROM4[194]<=16'd57245;
ROM1[195]<=16'd4712; ROM2[195]<=16'd0; ROM3[195]<=16'd23787; ROM4[195]<=16'd57245;
ROM1[196]<=16'd4673; ROM2[196]<=16'd0; ROM3[196]<=16'd23773; ROM4[196]<=16'd57225;
ROM1[197]<=16'd4662; ROM2[197]<=16'd0; ROM3[197]<=16'd23778; ROM4[197]<=16'd57222;
ROM1[198]<=16'd4688; ROM2[198]<=16'd0; ROM3[198]<=16'd23786; ROM4[198]<=16'd57234;
ROM1[199]<=16'd4729; ROM2[199]<=16'd0; ROM3[199]<=16'd23786; ROM4[199]<=16'd57245;
ROM1[200]<=16'd4749; ROM2[200]<=16'd0; ROM3[200]<=16'd23773; ROM4[200]<=16'd57244;
ROM1[201]<=16'd4734; ROM2[201]<=16'd0; ROM3[201]<=16'd23760; ROM4[201]<=16'd57232;
ROM1[202]<=16'd4713; ROM2[202]<=16'd0; ROM3[202]<=16'd23759; ROM4[202]<=16'd57228;
ROM1[203]<=16'd4692; ROM2[203]<=16'd0; ROM3[203]<=16'd23762; ROM4[203]<=16'd57224;
ROM1[204]<=16'd4682; ROM2[204]<=16'd0; ROM3[204]<=16'd23768; ROM4[204]<=16'd57224;
ROM1[205]<=16'd4677; ROM2[205]<=16'd0; ROM3[205]<=16'd23780; ROM4[205]<=16'd57233;
ROM1[206]<=16'd4679; ROM2[206]<=16'd0; ROM3[206]<=16'd23782; ROM4[206]<=16'd57235;
ROM1[207]<=16'd4696; ROM2[207]<=16'd0; ROM3[207]<=16'd23770; ROM4[207]<=16'd57233;
ROM1[208]<=16'd4727; ROM2[208]<=16'd0; ROM3[208]<=16'd23760; ROM4[208]<=16'd57235;
ROM1[209]<=16'd4735; ROM2[209]<=16'd0; ROM3[209]<=16'd23756; ROM4[209]<=16'd57233;
ROM1[210]<=16'd4723; ROM2[210]<=16'd0; ROM3[210]<=16'd23760; ROM4[210]<=16'd57233;
ROM1[211]<=16'd4704; ROM2[211]<=16'd0; ROM3[211]<=16'd23766; ROM4[211]<=16'd57230;
ROM1[212]<=16'd4694; ROM2[212]<=16'd0; ROM3[212]<=16'd23767; ROM4[212]<=16'd57230;
ROM1[213]<=16'd4681; ROM2[213]<=16'd0; ROM3[213]<=16'd23776; ROM4[213]<=16'd57234;
ROM1[214]<=16'd4671; ROM2[214]<=16'd0; ROM3[214]<=16'd23776; ROM4[214]<=16'd57235;
ROM1[215]<=16'd4685; ROM2[215]<=16'd0; ROM3[215]<=16'd23766; ROM4[215]<=16'd57232;
ROM1[216]<=16'd4730; ROM2[216]<=16'd0; ROM3[216]<=16'd23760; ROM4[216]<=16'd57236;
ROM1[217]<=16'd4770; ROM2[217]<=16'd0; ROM3[217]<=16'd23767; ROM4[217]<=16'd57257;
ROM1[218]<=16'd4759; ROM2[218]<=16'd0; ROM3[218]<=16'd23768; ROM4[218]<=16'd57256;
ROM1[219]<=16'd4735; ROM2[219]<=16'd0; ROM3[219]<=16'd23773; ROM4[219]<=16'd57250;
ROM1[220]<=16'd4715; ROM2[220]<=16'd0; ROM3[220]<=16'd23776; ROM4[220]<=16'd57247;
ROM1[221]<=16'd4687; ROM2[221]<=16'd0; ROM3[221]<=16'd23768; ROM4[221]<=16'd57233;
ROM1[222]<=16'd4692; ROM2[222]<=16'd0; ROM3[222]<=16'd23782; ROM4[222]<=16'd57239;
ROM1[223]<=16'd4717; ROM2[223]<=16'd0; ROM3[223]<=16'd23794; ROM4[223]<=16'd57254;
ROM1[224]<=16'd4737; ROM2[224]<=16'd0; ROM3[224]<=16'd23784; ROM4[224]<=16'd57249;
ROM1[225]<=16'd4755; ROM2[225]<=16'd0; ROM3[225]<=16'd23767; ROM4[225]<=16'd57241;
ROM1[226]<=16'd4758; ROM2[226]<=16'd0; ROM3[226]<=16'd23772; ROM4[226]<=16'd57246;
ROM1[227]<=16'd4741; ROM2[227]<=16'd0; ROM3[227]<=16'd23775; ROM4[227]<=16'd57245;
ROM1[228]<=16'd4734; ROM2[228]<=16'd0; ROM3[228]<=16'd23791; ROM4[228]<=16'd57255;
ROM1[229]<=16'd4727; ROM2[229]<=16'd0; ROM3[229]<=16'd23802; ROM4[229]<=16'd57263;
ROM1[230]<=16'd4689; ROM2[230]<=16'd0; ROM3[230]<=16'd23784; ROM4[230]<=16'd57242;
ROM1[231]<=16'd4682; ROM2[231]<=16'd0; ROM3[231]<=16'd23769; ROM4[231]<=16'd57230;
ROM1[232]<=16'd4698; ROM2[232]<=16'd0; ROM3[232]<=16'd23752; ROM4[232]<=16'd57224;
ROM1[233]<=16'd4728; ROM2[233]<=16'd0; ROM3[233]<=16'd23738; ROM4[233]<=16'd57220;
ROM1[234]<=16'd4746; ROM2[234]<=16'd0; ROM3[234]<=16'd23742; ROM4[234]<=16'd57228;
ROM1[235]<=16'd4736; ROM2[235]<=16'd0; ROM3[235]<=16'd23750; ROM4[235]<=16'd57231;
ROM1[236]<=16'd4714; ROM2[236]<=16'd0; ROM3[236]<=16'd23757; ROM4[236]<=16'd57230;
ROM1[237]<=16'd4697; ROM2[237]<=16'd0; ROM3[237]<=16'd23760; ROM4[237]<=16'd57230;
ROM1[238]<=16'd4689; ROM2[238]<=16'd0; ROM3[238]<=16'd23768; ROM4[238]<=16'd57235;
ROM1[239]<=16'd4691; ROM2[239]<=16'd0; ROM3[239]<=16'd23779; ROM4[239]<=16'd57243;
ROM1[240]<=16'd4697; ROM2[240]<=16'd0; ROM3[240]<=16'd23766; ROM4[240]<=16'd57234;
ROM1[241]<=16'd4733; ROM2[241]<=16'd0; ROM3[241]<=16'd23755; ROM4[241]<=16'd57236;
ROM1[242]<=16'd4761; ROM2[242]<=16'd0; ROM3[242]<=16'd23763; ROM4[242]<=16'd57246;
ROM1[243]<=16'd4723; ROM2[243]<=16'd0; ROM3[243]<=16'd23745; ROM4[243]<=16'd57224;
ROM1[244]<=16'd4688; ROM2[244]<=16'd0; ROM3[244]<=16'd23741; ROM4[244]<=16'd57213;
ROM1[245]<=16'd4681; ROM2[245]<=16'd0; ROM3[245]<=16'd23757; ROM4[245]<=16'd57222;
ROM1[246]<=16'd4657; ROM2[246]<=16'd0; ROM3[246]<=16'd23750; ROM4[246]<=16'd57215;
ROM1[247]<=16'd4665; ROM2[247]<=16'd0; ROM3[247]<=16'd23763; ROM4[247]<=16'd57226;
ROM1[248]<=16'd4690; ROM2[248]<=16'd0; ROM3[248]<=16'd23774; ROM4[248]<=16'd57238;
ROM1[249]<=16'd4703; ROM2[249]<=16'd0; ROM3[249]<=16'd23759; ROM4[249]<=16'd57228;
ROM1[250]<=16'd4730; ROM2[250]<=16'd0; ROM3[250]<=16'd23752; ROM4[250]<=16'd57225;
ROM1[251]<=16'd4721; ROM2[251]<=16'd0; ROM3[251]<=16'd23748; ROM4[251]<=16'd57223;
ROM1[252]<=16'd4701; ROM2[252]<=16'd0; ROM3[252]<=16'd23750; ROM4[252]<=16'd57224;
ROM1[253]<=16'd4692; ROM2[253]<=16'd0; ROM3[253]<=16'd23761; ROM4[253]<=16'd57225;
ROM1[254]<=16'd4671; ROM2[254]<=16'd0; ROM3[254]<=16'd23756; ROM4[254]<=16'd57218;
ROM1[255]<=16'd4655; ROM2[255]<=16'd0; ROM3[255]<=16'd23757; ROM4[255]<=16'd57217;
ROM1[256]<=16'd4660; ROM2[256]<=16'd0; ROM3[256]<=16'd23760; ROM4[256]<=16'd57221;
ROM1[257]<=16'd4674; ROM2[257]<=16'd0; ROM3[257]<=16'd23742; ROM4[257]<=16'd57217;
ROM1[258]<=16'd4703; ROM2[258]<=16'd0; ROM3[258]<=16'd23724; ROM4[258]<=16'd57208;
ROM1[259]<=16'd4720; ROM2[259]<=16'd0; ROM3[259]<=16'd23725; ROM4[259]<=16'd57210;
ROM1[260]<=16'd4706; ROM2[260]<=16'd0; ROM3[260]<=16'd23729; ROM4[260]<=16'd57210;
ROM1[261]<=16'd4688; ROM2[261]<=16'd0; ROM3[261]<=16'd23739; ROM4[261]<=16'd57212;
ROM1[262]<=16'd4670; ROM2[262]<=16'd0; ROM3[262]<=16'd23746; ROM4[262]<=16'd57214;
ROM1[263]<=16'd4648; ROM2[263]<=16'd0; ROM3[263]<=16'd23750; ROM4[263]<=16'd57209;
ROM1[264]<=16'd4650; ROM2[264]<=16'd0; ROM3[264]<=16'd23761; ROM4[264]<=16'd57215;
ROM1[265]<=16'd4674; ROM2[265]<=16'd0; ROM3[265]<=16'd23764; ROM4[265]<=16'd57223;
ROM1[266]<=16'd4716; ROM2[266]<=16'd0; ROM3[266]<=16'd23763; ROM4[266]<=16'd57233;
ROM1[267]<=16'd4752; ROM2[267]<=16'd0; ROM3[267]<=16'd23772; ROM4[267]<=16'd57252;
ROM1[268]<=16'd4754; ROM2[268]<=16'd0; ROM3[268]<=16'd23784; ROM4[268]<=16'd57261;
ROM1[269]<=16'd4729; ROM2[269]<=16'd0; ROM3[269]<=16'd23780; ROM4[269]<=16'd57255;
ROM1[270]<=16'd4709; ROM2[270]<=16'd0; ROM3[270]<=16'd23779; ROM4[270]<=16'd57249;
ROM1[271]<=16'd4690; ROM2[271]<=16'd0; ROM3[271]<=16'd23785; ROM4[271]<=16'd57244;
ROM1[272]<=16'd4675; ROM2[272]<=16'd0; ROM3[272]<=16'd23778; ROM4[272]<=16'd57238;
ROM1[273]<=16'd4687; ROM2[273]<=16'd0; ROM3[273]<=16'd23778; ROM4[273]<=16'd57239;
ROM1[274]<=16'd4718; ROM2[274]<=16'd0; ROM3[274]<=16'd23773; ROM4[274]<=16'd57244;
ROM1[275]<=16'd4735; ROM2[275]<=16'd0; ROM3[275]<=16'd23749; ROM4[275]<=16'd57233;
ROM1[276]<=16'd4727; ROM2[276]<=16'd0; ROM3[276]<=16'd23745; ROM4[276]<=16'd57228;
ROM1[277]<=16'd4722; ROM2[277]<=16'd0; ROM3[277]<=16'd23762; ROM4[277]<=16'd57235;
ROM1[278]<=16'd4709; ROM2[278]<=16'd0; ROM3[278]<=16'd23773; ROM4[278]<=16'd57239;
ROM1[279]<=16'd4714; ROM2[279]<=16'd0; ROM3[279]<=16'd23790; ROM4[279]<=16'd57253;
ROM1[280]<=16'd4705; ROM2[280]<=16'd0; ROM3[280]<=16'd23793; ROM4[280]<=16'd57250;
ROM1[281]<=16'd4690; ROM2[281]<=16'd0; ROM3[281]<=16'd23781; ROM4[281]<=16'd57237;
ROM1[282]<=16'd4710; ROM2[282]<=16'd0; ROM3[282]<=16'd23771; ROM4[282]<=16'd57234;
ROM1[283]<=16'd4729; ROM2[283]<=16'd0; ROM3[283]<=16'd23752; ROM4[283]<=16'd57225;
ROM1[284]<=16'd4722; ROM2[284]<=16'd0; ROM3[284]<=16'd23746; ROM4[284]<=16'd57222;
ROM1[285]<=16'd4706; ROM2[285]<=16'd0; ROM3[285]<=16'd23749; ROM4[285]<=16'd57219;
ROM1[286]<=16'd4696; ROM2[286]<=16'd0; ROM3[286]<=16'd23763; ROM4[286]<=16'd57230;
ROM1[287]<=16'd4692; ROM2[287]<=16'd0; ROM3[287]<=16'd23781; ROM4[287]<=16'd57242;
ROM1[288]<=16'd4677; ROM2[288]<=16'd0; ROM3[288]<=16'd23781; ROM4[288]<=16'd57238;
ROM1[289]<=16'd4662; ROM2[289]<=16'd0; ROM3[289]<=16'd23769; ROM4[289]<=16'd57225;
ROM1[290]<=16'd4669; ROM2[290]<=16'd0; ROM3[290]<=16'd23756; ROM4[290]<=16'd57217;
ROM1[291]<=16'd4698; ROM2[291]<=16'd0; ROM3[291]<=16'd23745; ROM4[291]<=16'd57218;
ROM1[292]<=16'd4727; ROM2[292]<=16'd0; ROM3[292]<=16'd23745; ROM4[292]<=16'd57229;
ROM1[293]<=16'd4732; ROM2[293]<=16'd0; ROM3[293]<=16'd23763; ROM4[293]<=16'd57241;
ROM1[294]<=16'd4722; ROM2[294]<=16'd0; ROM3[294]<=16'd23783; ROM4[294]<=16'd57250;
ROM1[295]<=16'd4708; ROM2[295]<=16'd0; ROM3[295]<=16'd23789; ROM4[295]<=16'd57250;
ROM1[296]<=16'd4694; ROM2[296]<=16'd0; ROM3[296]<=16'd23792; ROM4[296]<=16'd57254;
ROM1[297]<=16'd4670; ROM2[297]<=16'd0; ROM3[297]<=16'd23777; ROM4[297]<=16'd57235;
ROM1[298]<=16'd4658; ROM2[298]<=16'd0; ROM3[298]<=16'd23751; ROM4[298]<=16'd57213;
ROM1[299]<=16'd4684; ROM2[299]<=16'd0; ROM3[299]<=16'd23738; ROM4[299]<=16'd57213;
ROM1[300]<=16'd4704; ROM2[300]<=16'd0; ROM3[300]<=16'd23726; ROM4[300]<=16'd57210;
ROM1[301]<=16'd4705; ROM2[301]<=16'd0; ROM3[301]<=16'd23733; ROM4[301]<=16'd57220;
ROM1[302]<=16'd4684; ROM2[302]<=16'd0; ROM3[302]<=16'd23738; ROM4[302]<=16'd57218;
ROM1[303]<=16'd4662; ROM2[303]<=16'd0; ROM3[303]<=16'd23744; ROM4[303]<=16'd57215;
ROM1[304]<=16'd4662; ROM2[304]<=16'd0; ROM3[304]<=16'd23760; ROM4[304]<=16'd57221;
ROM1[305]<=16'd4665; ROM2[305]<=16'd0; ROM3[305]<=16'd23776; ROM4[305]<=16'd57232;
ROM1[306]<=16'd4673; ROM2[306]<=16'd0; ROM3[306]<=16'd23784; ROM4[306]<=16'd57239;
ROM1[307]<=16'd4687; ROM2[307]<=16'd0; ROM3[307]<=16'd23767; ROM4[307]<=16'd57228;
ROM1[308]<=16'd4716; ROM2[308]<=16'd0; ROM3[308]<=16'd23746; ROM4[308]<=16'd57221;
ROM1[309]<=16'd4718; ROM2[309]<=16'd0; ROM3[309]<=16'd23738; ROM4[309]<=16'd57217;
ROM1[310]<=16'd4702; ROM2[310]<=16'd0; ROM3[310]<=16'd23744; ROM4[310]<=16'd57220;
ROM1[311]<=16'd4696; ROM2[311]<=16'd0; ROM3[311]<=16'd23761; ROM4[311]<=16'd57229;
ROM1[312]<=16'd4695; ROM2[312]<=16'd0; ROM3[312]<=16'd23778; ROM4[312]<=16'd57240;
ROM1[313]<=16'd4698; ROM2[313]<=16'd0; ROM3[313]<=16'd23802; ROM4[313]<=16'd57258;
ROM1[314]<=16'd4704; ROM2[314]<=16'd0; ROM3[314]<=16'd23804; ROM4[314]<=16'd57259;
ROM1[315]<=16'd4702; ROM2[315]<=16'd0; ROM3[315]<=16'd23784; ROM4[315]<=16'd57242;
ROM1[316]<=16'd4730; ROM2[316]<=16'd0; ROM3[316]<=16'd23773; ROM4[316]<=16'd57240;
ROM1[317]<=16'd4751; ROM2[317]<=16'd0; ROM3[317]<=16'd23759; ROM4[317]<=16'd57237;
ROM1[318]<=16'd4733; ROM2[318]<=16'd0; ROM3[318]<=16'd23751; ROM4[318]<=16'd57230;
ROM1[319]<=16'd4714; ROM2[319]<=16'd0; ROM3[319]<=16'd23760; ROM4[319]<=16'd57229;
ROM1[320]<=16'd4702; ROM2[320]<=16'd0; ROM3[320]<=16'd23770; ROM4[320]<=16'd57238;
ROM1[321]<=16'd4681; ROM2[321]<=16'd0; ROM3[321]<=16'd23769; ROM4[321]<=16'd57236;
ROM1[322]<=16'd4673; ROM2[322]<=16'd0; ROM3[322]<=16'd23772; ROM4[322]<=16'd57238;
ROM1[323]<=16'd4692; ROM2[323]<=16'd0; ROM3[323]<=16'd23776; ROM4[323]<=16'd57247;
ROM1[324]<=16'd4712; ROM2[324]<=16'd0; ROM3[324]<=16'd23759; ROM4[324]<=16'd57238;
ROM1[325]<=16'd4744; ROM2[325]<=16'd0; ROM3[325]<=16'd23754; ROM4[325]<=16'd57242;
ROM1[326]<=16'd4759; ROM2[326]<=16'd0; ROM3[326]<=16'd23769; ROM4[326]<=16'd57257;
ROM1[327]<=16'd4749; ROM2[327]<=16'd0; ROM3[327]<=16'd23785; ROM4[327]<=16'd57264;
ROM1[328]<=16'd4713; ROM2[328]<=16'd0; ROM3[328]<=16'd23780; ROM4[328]<=16'd57246;
ROM1[329]<=16'd4676; ROM2[329]<=16'd0; ROM3[329]<=16'd23769; ROM4[329]<=16'd57226;
ROM1[330]<=16'd4656; ROM2[330]<=16'd0; ROM3[330]<=16'd23772; ROM4[330]<=16'd57224;
ROM1[331]<=16'd4667; ROM2[331]<=16'd0; ROM3[331]<=16'd23777; ROM4[331]<=16'd57228;
ROM1[332]<=16'd4706; ROM2[332]<=16'd0; ROM3[332]<=16'd23781; ROM4[332]<=16'd57239;
ROM1[333]<=16'd4746; ROM2[333]<=16'd0; ROM3[333]<=16'd23781; ROM4[333]<=16'd57251;
ROM1[334]<=16'd4761; ROM2[334]<=16'd0; ROM3[334]<=16'd23787; ROM4[334]<=16'd57254;
ROM1[335]<=16'd4730; ROM2[335]<=16'd0; ROM3[335]<=16'd23776; ROM4[335]<=16'd57241;
ROM1[336]<=16'd4698; ROM2[336]<=16'd0; ROM3[336]<=16'd23772; ROM4[336]<=16'd57235;
ROM1[337]<=16'd4689; ROM2[337]<=16'd0; ROM3[337]<=16'd23781; ROM4[337]<=16'd57237;
ROM1[338]<=16'd4674; ROM2[338]<=16'd0; ROM3[338]<=16'd23781; ROM4[338]<=16'd57232;
ROM1[339]<=16'd4671; ROM2[339]<=16'd0; ROM3[339]<=16'd23788; ROM4[339]<=16'd57236;
ROM1[340]<=16'd4691; ROM2[340]<=16'd0; ROM3[340]<=16'd23788; ROM4[340]<=16'd57238;
ROM1[341]<=16'd4720; ROM2[341]<=16'd0; ROM3[341]<=16'd23768; ROM4[341]<=16'd57234;
ROM1[342]<=16'd4723; ROM2[342]<=16'd0; ROM3[342]<=16'd23745; ROM4[342]<=16'd57220;
ROM1[343]<=16'd4712; ROM2[343]<=16'd0; ROM3[343]<=16'd23742; ROM4[343]<=16'd57213;
ROM1[344]<=16'd4699; ROM2[344]<=16'd0; ROM3[344]<=16'd23751; ROM4[344]<=16'd57218;
ROM1[345]<=16'd4683; ROM2[345]<=16'd0; ROM3[345]<=16'd23757; ROM4[345]<=16'd57219;
ROM1[346]<=16'd4671; ROM2[346]<=16'd0; ROM3[346]<=16'd23767; ROM4[346]<=16'd57224;
ROM1[347]<=16'd4670; ROM2[347]<=16'd0; ROM3[347]<=16'd23775; ROM4[347]<=16'd57231;
ROM1[348]<=16'd4677; ROM2[348]<=16'd0; ROM3[348]<=16'd23767; ROM4[348]<=16'd57226;
ROM1[349]<=16'd4702; ROM2[349]<=16'd0; ROM3[349]<=16'd23756; ROM4[349]<=16'd57225;
ROM1[350]<=16'd4733; ROM2[350]<=16'd0; ROM3[350]<=16'd23750; ROM4[350]<=16'd57232;
ROM1[351]<=16'd4737; ROM2[351]<=16'd0; ROM3[351]<=16'd23759; ROM4[351]<=16'd57239;
ROM1[352]<=16'd4728; ROM2[352]<=16'd0; ROM3[352]<=16'd23777; ROM4[352]<=16'd57248;
ROM1[353]<=16'd4707; ROM2[353]<=16'd0; ROM3[353]<=16'd23785; ROM4[353]<=16'd57245;
ROM1[354]<=16'd4692; ROM2[354]<=16'd0; ROM3[354]<=16'd23788; ROM4[354]<=16'd57243;
ROM1[355]<=16'd4678; ROM2[355]<=16'd0; ROM3[355]<=16'd23788; ROM4[355]<=16'd57239;
ROM1[356]<=16'd4678; ROM2[356]<=16'd0; ROM3[356]<=16'd23785; ROM4[356]<=16'd57235;
ROM1[357]<=16'd4699; ROM2[357]<=16'd0; ROM3[357]<=16'd23777; ROM4[357]<=16'd57239;
ROM1[358]<=16'd4731; ROM2[358]<=16'd0; ROM3[358]<=16'd23764; ROM4[358]<=16'd57243;
ROM1[359]<=16'd4730; ROM2[359]<=16'd0; ROM3[359]<=16'd23754; ROM4[359]<=16'd57236;
ROM1[360]<=16'd4710; ROM2[360]<=16'd0; ROM3[360]<=16'd23754; ROM4[360]<=16'd57232;
ROM1[361]<=16'd4705; ROM2[361]<=16'd0; ROM3[361]<=16'd23774; ROM4[361]<=16'd57244;
ROM1[362]<=16'd4713; ROM2[362]<=16'd0; ROM3[362]<=16'd23800; ROM4[362]<=16'd57263;
ROM1[363]<=16'd4684; ROM2[363]<=16'd0; ROM3[363]<=16'd23792; ROM4[363]<=16'd57256;
ROM1[364]<=16'd4669; ROM2[364]<=16'd0; ROM3[364]<=16'd23783; ROM4[364]<=16'd57246;
ROM1[365]<=16'd4691; ROM2[365]<=16'd0; ROM3[365]<=16'd23779; ROM4[365]<=16'd57245;
ROM1[366]<=16'd4717; ROM2[366]<=16'd0; ROM3[366]<=16'd23758; ROM4[366]<=16'd57235;
ROM1[367]<=16'd4755; ROM2[367]<=16'd0; ROM3[367]<=16'd23766; ROM4[367]<=16'd57250;
ROM1[368]<=16'd4768; ROM2[368]<=16'd0; ROM3[368]<=16'd23788; ROM4[368]<=16'd57269;
ROM1[369]<=16'd4744; ROM2[369]<=16'd0; ROM3[369]<=16'd23791; ROM4[369]<=16'd57266;
ROM1[370]<=16'd4717; ROM2[370]<=16'd0; ROM3[370]<=16'd23792; ROM4[370]<=16'd57258;
ROM1[371]<=16'd4686; ROM2[371]<=16'd0; ROM3[371]<=16'd23786; ROM4[371]<=16'd57244;
ROM1[372]<=16'd4678; ROM2[372]<=16'd0; ROM3[372]<=16'd23782; ROM4[372]<=16'd57239;
ROM1[373]<=16'd4690; ROM2[373]<=16'd0; ROM3[373]<=16'd23775; ROM4[373]<=16'd57232;
ROM1[374]<=16'd4713; ROM2[374]<=16'd0; ROM3[374]<=16'd23763; ROM4[374]<=16'd57230;
ROM1[375]<=16'd4746; ROM2[375]<=16'd0; ROM3[375]<=16'd23768; ROM4[375]<=16'd57242;
ROM1[376]<=16'd4742; ROM2[376]<=16'd0; ROM3[376]<=16'd23776; ROM4[376]<=16'd57246;
ROM1[377]<=16'd4720; ROM2[377]<=16'd0; ROM3[377]<=16'd23779; ROM4[377]<=16'd57241;
ROM1[378]<=16'd4705; ROM2[378]<=16'd0; ROM3[378]<=16'd23782; ROM4[378]<=16'd57237;
ROM1[379]<=16'd4692; ROM2[379]<=16'd0; ROM3[379]<=16'd23786; ROM4[379]<=16'd57238;
ROM1[380]<=16'd4684; ROM2[380]<=16'd0; ROM3[380]<=16'd23793; ROM4[380]<=16'd57242;
ROM1[381]<=16'd4695; ROM2[381]<=16'd0; ROM3[381]<=16'd23805; ROM4[381]<=16'd57253;
ROM1[382]<=16'd4736; ROM2[382]<=16'd0; ROM3[382]<=16'd23818; ROM4[382]<=16'd57273;
ROM1[383]<=16'd4771; ROM2[383]<=16'd0; ROM3[383]<=16'd23804; ROM4[383]<=16'd57272;
ROM1[384]<=16'd4750; ROM2[384]<=16'd0; ROM3[384]<=16'd23769; ROM4[384]<=16'd57242;
ROM1[385]<=16'd4721; ROM2[385]<=16'd0; ROM3[385]<=16'd23763; ROM4[385]<=16'd57231;
ROM1[386]<=16'd4705; ROM2[386]<=16'd0; ROM3[386]<=16'd23774; ROM4[386]<=16'd57234;
ROM1[387]<=16'd4693; ROM2[387]<=16'd0; ROM3[387]<=16'd23780; ROM4[387]<=16'd57230;
ROM1[388]<=16'd4679; ROM2[388]<=16'd0; ROM3[388]<=16'd23787; ROM4[388]<=16'd57233;
ROM1[389]<=16'd4674; ROM2[389]<=16'd0; ROM3[389]<=16'd23781; ROM4[389]<=16'd57227;
ROM1[390]<=16'd4676; ROM2[390]<=16'd0; ROM3[390]<=16'd23764; ROM4[390]<=16'd57210;
ROM1[391]<=16'd4711; ROM2[391]<=16'd0; ROM3[391]<=16'd23753; ROM4[391]<=16'd57211;
ROM1[392]<=16'd4743; ROM2[392]<=16'd0; ROM3[392]<=16'd23757; ROM4[392]<=16'd57225;
ROM1[393]<=16'd4731; ROM2[393]<=16'd0; ROM3[393]<=16'd23760; ROM4[393]<=16'd57225;
ROM1[394]<=16'd4705; ROM2[394]<=16'd0; ROM3[394]<=16'd23756; ROM4[394]<=16'd57215;
ROM1[395]<=16'd4693; ROM2[395]<=16'd0; ROM3[395]<=16'd23765; ROM4[395]<=16'd57218;
ROM1[396]<=16'd4682; ROM2[396]<=16'd0; ROM3[396]<=16'd23772; ROM4[396]<=16'd57220;
ROM1[397]<=16'd4677; ROM2[397]<=16'd0; ROM3[397]<=16'd23774; ROM4[397]<=16'd57218;
ROM1[398]<=16'd4694; ROM2[398]<=16'd0; ROM3[398]<=16'd23780; ROM4[398]<=16'd57230;
ROM1[399]<=16'd4723; ROM2[399]<=16'd0; ROM3[399]<=16'd23769; ROM4[399]<=16'd57231;
ROM1[400]<=16'd4748; ROM2[400]<=16'd0; ROM3[400]<=16'd23751; ROM4[400]<=16'd57226;
ROM1[401]<=16'd4739; ROM2[401]<=16'd0; ROM3[401]<=16'd23747; ROM4[401]<=16'd57221;
ROM1[402]<=16'd4714; ROM2[402]<=16'd0; ROM3[402]<=16'd23746; ROM4[402]<=16'd57215;
ROM1[403]<=16'd4698; ROM2[403]<=16'd0; ROM3[403]<=16'd23757; ROM4[403]<=16'd57218;
ROM1[404]<=16'd4684; ROM2[404]<=16'd0; ROM3[404]<=16'd23776; ROM4[404]<=16'd57227;
ROM1[405]<=16'd4677; ROM2[405]<=16'd0; ROM3[405]<=16'd23786; ROM4[405]<=16'd57235;
ROM1[406]<=16'd4686; ROM2[406]<=16'd0; ROM3[406]<=16'd23786; ROM4[406]<=16'd57237;
ROM1[407]<=16'd4707; ROM2[407]<=16'd0; ROM3[407]<=16'd23781; ROM4[407]<=16'd57240;
ROM1[408]<=16'd4740; ROM2[408]<=16'd0; ROM3[408]<=16'd23770; ROM4[408]<=16'd57240;
ROM1[409]<=16'd4769; ROM2[409]<=16'd0; ROM3[409]<=16'd23787; ROM4[409]<=16'd57260;
ROM1[410]<=16'd4767; ROM2[410]<=16'd0; ROM3[410]<=16'd23806; ROM4[410]<=16'd57273;
ROM1[411]<=16'd4732; ROM2[411]<=16'd0; ROM3[411]<=16'd23797; ROM4[411]<=16'd57256;
ROM1[412]<=16'd4727; ROM2[412]<=16'd0; ROM3[412]<=16'd23808; ROM4[412]<=16'd57265;
ROM1[413]<=16'd4710; ROM2[413]<=16'd0; ROM3[413]<=16'd23813; ROM4[413]<=16'd57265;
ROM1[414]<=16'd4701; ROM2[414]<=16'd0; ROM3[414]<=16'd23809; ROM4[414]<=16'd57261;
ROM1[415]<=16'd4729; ROM2[415]<=16'd0; ROM3[415]<=16'd23811; ROM4[415]<=16'd57270;
ROM1[416]<=16'd4762; ROM2[416]<=16'd0; ROM3[416]<=16'd23798; ROM4[416]<=16'd57265;
ROM1[417]<=16'd4774; ROM2[417]<=16'd0; ROM3[417]<=16'd23787; ROM4[417]<=16'd57264;
ROM1[418]<=16'd4770; ROM2[418]<=16'd0; ROM3[418]<=16'd23803; ROM4[418]<=16'd57276;
ROM1[419]<=16'd4754; ROM2[419]<=16'd0; ROM3[419]<=16'd23816; ROM4[419]<=16'd57280;
ROM1[420]<=16'd4727; ROM2[420]<=16'd0; ROM3[420]<=16'd23810; ROM4[420]<=16'd57269;
ROM1[421]<=16'd4706; ROM2[421]<=16'd0; ROM3[421]<=16'd23807; ROM4[421]<=16'd57259;
ROM1[422]<=16'd4691; ROM2[422]<=16'd0; ROM3[422]<=16'd23797; ROM4[422]<=16'd57247;
ROM1[423]<=16'd4707; ROM2[423]<=16'd0; ROM3[423]<=16'd23798; ROM4[423]<=16'd57252;
ROM1[424]<=16'd4737; ROM2[424]<=16'd0; ROM3[424]<=16'd23795; ROM4[424]<=16'd57260;
ROM1[425]<=16'd4749; ROM2[425]<=16'd0; ROM3[425]<=16'd23777; ROM4[425]<=16'd57252;
ROM1[426]<=16'd4745; ROM2[426]<=16'd0; ROM3[426]<=16'd23775; ROM4[426]<=16'd57249;
ROM1[427]<=16'd4729; ROM2[427]<=16'd0; ROM3[427]<=16'd23786; ROM4[427]<=16'd57251;
ROM1[428]<=16'd4714; ROM2[428]<=16'd0; ROM3[428]<=16'd23798; ROM4[428]<=16'd57254;
ROM1[429]<=16'd4711; ROM2[429]<=16'd0; ROM3[429]<=16'd23812; ROM4[429]<=16'd57264;
ROM1[430]<=16'd4710; ROM2[430]<=16'd0; ROM3[430]<=16'd23824; ROM4[430]<=16'd57272;
ROM1[431]<=16'd4715; ROM2[431]<=16'd0; ROM3[431]<=16'd23828; ROM4[431]<=16'd57275;
ROM1[432]<=16'd4745; ROM2[432]<=16'd0; ROM3[432]<=16'd23830; ROM4[432]<=16'd57281;
ROM1[433]<=16'd4779; ROM2[433]<=16'd0; ROM3[433]<=16'd23822; ROM4[433]<=16'd57282;
ROM1[434]<=16'd4752; ROM2[434]<=16'd0; ROM3[434]<=16'd23788; ROM4[434]<=16'd57253;
ROM1[435]<=16'd4715; ROM2[435]<=16'd0; ROM3[435]<=16'd23772; ROM4[435]<=16'd57235;
ROM1[436]<=16'd4703; ROM2[436]<=16'd0; ROM3[436]<=16'd23782; ROM4[436]<=16'd57239;
ROM1[437]<=16'd4699; ROM2[437]<=16'd0; ROM3[437]<=16'd23791; ROM4[437]<=16'd57243;
ROM1[438]<=16'd4697; ROM2[438]<=16'd0; ROM3[438]<=16'd23810; ROM4[438]<=16'd57256;
ROM1[439]<=16'd4702; ROM2[439]<=16'd0; ROM3[439]<=16'd23816; ROM4[439]<=16'd57261;
ROM1[440]<=16'd4729; ROM2[440]<=16'd0; ROM3[440]<=16'd23816; ROM4[440]<=16'd57266;
ROM1[441]<=16'd4776; ROM2[441]<=16'd0; ROM3[441]<=16'd23823; ROM4[441]<=16'd57286;
ROM1[442]<=16'd4800; ROM2[442]<=16'd0; ROM3[442]<=16'd23828; ROM4[442]<=16'd57293;
ROM1[443]<=16'd4779; ROM2[443]<=16'd0; ROM3[443]<=16'd23823; ROM4[443]<=16'd57284;
ROM1[444]<=16'd4744; ROM2[444]<=16'd0; ROM3[444]<=16'd23814; ROM4[444]<=16'd57265;
ROM1[445]<=16'd4720; ROM2[445]<=16'd0; ROM3[445]<=16'd23804; ROM4[445]<=16'd57253;
ROM1[446]<=16'd4703; ROM2[446]<=16'd0; ROM3[446]<=16'd23805; ROM4[446]<=16'd57249;
ROM1[447]<=16'd4703; ROM2[447]<=16'd0; ROM3[447]<=16'd23821; ROM4[447]<=16'd57256;
ROM1[448]<=16'd4703; ROM2[448]<=16'd0; ROM3[448]<=16'd23815; ROM4[448]<=16'd57255;
ROM1[449]<=16'd4723; ROM2[449]<=16'd0; ROM3[449]<=16'd23797; ROM4[449]<=16'd57247;
ROM1[450]<=16'd4753; ROM2[450]<=16'd0; ROM3[450]<=16'd23786; ROM4[450]<=16'd57246;
ROM1[451]<=16'd4747; ROM2[451]<=16'd0; ROM3[451]<=16'd23781; ROM4[451]<=16'd57243;
ROM1[452]<=16'd4738; ROM2[452]<=16'd0; ROM3[452]<=16'd23794; ROM4[452]<=16'd57251;
ROM1[453]<=16'd4732; ROM2[453]<=16'd0; ROM3[453]<=16'd23808; ROM4[453]<=16'd57256;
ROM1[454]<=16'd4717; ROM2[454]<=16'd0; ROM3[454]<=16'd23809; ROM4[454]<=16'd57252;
ROM1[455]<=16'd4706; ROM2[455]<=16'd0; ROM3[455]<=16'd23816; ROM4[455]<=16'd57251;
ROM1[456]<=16'd4709; ROM2[456]<=16'd0; ROM3[456]<=16'd23812; ROM4[456]<=16'd57247;
ROM1[457]<=16'd4722; ROM2[457]<=16'd0; ROM3[457]<=16'd23791; ROM4[457]<=16'd57238;
ROM1[458]<=16'd4756; ROM2[458]<=16'd0; ROM3[458]<=16'd23782; ROM4[458]<=16'd57242;
ROM1[459]<=16'd4770; ROM2[459]<=16'd0; ROM3[459]<=16'd23783; ROM4[459]<=16'd57252;
ROM1[460]<=16'd4753; ROM2[460]<=16'd0; ROM3[460]<=16'd23790; ROM4[460]<=16'd57255;
ROM1[461]<=16'd4735; ROM2[461]<=16'd0; ROM3[461]<=16'd23799; ROM4[461]<=16'd57254;
ROM1[462]<=16'd4717; ROM2[462]<=16'd0; ROM3[462]<=16'd23800; ROM4[462]<=16'd57249;
ROM1[463]<=16'd4704; ROM2[463]<=16'd0; ROM3[463]<=16'd23808; ROM4[463]<=16'd57249;
ROM1[464]<=16'd4702; ROM2[464]<=16'd0; ROM3[464]<=16'd23812; ROM4[464]<=16'd57252;
ROM1[465]<=16'd4710; ROM2[465]<=16'd0; ROM3[465]<=16'd23801; ROM4[465]<=16'd57251;
ROM1[466]<=16'd4744; ROM2[466]<=16'd0; ROM3[466]<=16'd23795; ROM4[466]<=16'd57256;
ROM1[467]<=16'd4768; ROM2[467]<=16'd0; ROM3[467]<=16'd23793; ROM4[467]<=16'd57259;
ROM1[468]<=16'd4749; ROM2[468]<=16'd0; ROM3[468]<=16'd23782; ROM4[468]<=16'd57246;
ROM1[469]<=16'd4739; ROM2[469]<=16'd0; ROM3[469]<=16'd23795; ROM4[469]<=16'd57250;
ROM1[470]<=16'd4735; ROM2[470]<=16'd0; ROM3[470]<=16'd23807; ROM4[470]<=16'd57257;
ROM1[471]<=16'd4716; ROM2[471]<=16'd0; ROM3[471]<=16'd23804; ROM4[471]<=16'd57256;
ROM1[472]<=16'd4707; ROM2[472]<=16'd0; ROM3[472]<=16'd23806; ROM4[472]<=16'd57255;
ROM1[473]<=16'd4707; ROM2[473]<=16'd0; ROM3[473]<=16'd23801; ROM4[473]<=16'd57248;
ROM1[474]<=16'd4729; ROM2[474]<=16'd0; ROM3[474]<=16'd23793; ROM4[474]<=16'd57239;
ROM1[475]<=16'd4754; ROM2[475]<=16'd0; ROM3[475]<=16'd23784; ROM4[475]<=16'd57237;
ROM1[476]<=16'd4760; ROM2[476]<=16'd0; ROM3[476]<=16'd23795; ROM4[476]<=16'd57244;
ROM1[477]<=16'd4758; ROM2[477]<=16'd0; ROM3[477]<=16'd23820; ROM4[477]<=16'd57263;
ROM1[478]<=16'd4732; ROM2[478]<=16'd0; ROM3[478]<=16'd23822; ROM4[478]<=16'd57260;
ROM1[479]<=16'd4702; ROM2[479]<=16'd0; ROM3[479]<=16'd23815; ROM4[479]<=16'd57245;
ROM1[480]<=16'd4703; ROM2[480]<=16'd0; ROM3[480]<=16'd23832; ROM4[480]<=16'd57257;
ROM1[481]<=16'd4728; ROM2[481]<=16'd0; ROM3[481]<=16'd23851; ROM4[481]<=16'd57275;
ROM1[482]<=16'd4737; ROM2[482]<=16'd0; ROM3[482]<=16'd23825; ROM4[482]<=16'd57260;
ROM1[483]<=16'd4756; ROM2[483]<=16'd0; ROM3[483]<=16'd23799; ROM4[483]<=16'd57249;
ROM1[484]<=16'd4751; ROM2[484]<=16'd0; ROM3[484]<=16'd23785; ROM4[484]<=16'd57239;
ROM1[485]<=16'd4718; ROM2[485]<=16'd0; ROM3[485]<=16'd23769; ROM4[485]<=16'd57221;
ROM1[486]<=16'd4706; ROM2[486]<=16'd0; ROM3[486]<=16'd23780; ROM4[486]<=16'd57227;
ROM1[487]<=16'd4705; ROM2[487]<=16'd0; ROM3[487]<=16'd23798; ROM4[487]<=16'd57237;
ROM1[488]<=16'd4690; ROM2[488]<=16'd0; ROM3[488]<=16'd23803; ROM4[488]<=16'd57239;
ROM1[489]<=16'd4688; ROM2[489]<=16'd0; ROM3[489]<=16'd23797; ROM4[489]<=16'd57234;
ROM1[490]<=16'd4710; ROM2[490]<=16'd0; ROM3[490]<=16'd23796; ROM4[490]<=16'd57240;
ROM1[491]<=16'd4738; ROM2[491]<=16'd0; ROM3[491]<=16'd23784; ROM4[491]<=16'd57242;
ROM1[492]<=16'd4752; ROM2[492]<=16'd0; ROM3[492]<=16'd23774; ROM4[492]<=16'd57239;
ROM1[493]<=16'd4736; ROM2[493]<=16'd0; ROM3[493]<=16'd23773; ROM4[493]<=16'd57238;
ROM1[494]<=16'd4717; ROM2[494]<=16'd0; ROM3[494]<=16'd23781; ROM4[494]<=16'd57241;
ROM1[495]<=16'd4705; ROM2[495]<=16'd0; ROM3[495]<=16'd23791; ROM4[495]<=16'd57243;
ROM1[496]<=16'd4696; ROM2[496]<=16'd0; ROM3[496]<=16'd23800; ROM4[496]<=16'd57250;
ROM1[497]<=16'd4691; ROM2[497]<=16'd0; ROM3[497]<=16'd23811; ROM4[497]<=16'd57256;
ROM1[498]<=16'd4702; ROM2[498]<=16'd0; ROM3[498]<=16'd23808; ROM4[498]<=16'd57254;
ROM1[499]<=16'd4736; ROM2[499]<=16'd0; ROM3[499]<=16'd23803; ROM4[499]<=16'd57260;
ROM1[500]<=16'd4772; ROM2[500]<=16'd0; ROM3[500]<=16'd23798; ROM4[500]<=16'd57268;
ROM1[501]<=16'd4771; ROM2[501]<=16'd0; ROM3[501]<=16'd23804; ROM4[501]<=16'd57268;
ROM1[502]<=16'd4752; ROM2[502]<=16'd0; ROM3[502]<=16'd23807; ROM4[502]<=16'd57264;
ROM1[503]<=16'd4733; ROM2[503]<=16'd0; ROM3[503]<=16'd23806; ROM4[503]<=16'd57259;
ROM1[504]<=16'd4719; ROM2[504]<=16'd0; ROM3[504]<=16'd23811; ROM4[504]<=16'd57258;
ROM1[505]<=16'd4696; ROM2[505]<=16'd0; ROM3[505]<=16'd23803; ROM4[505]<=16'd57249;
ROM1[506]<=16'd4695; ROM2[506]<=16'd0; ROM3[506]<=16'd23797; ROM4[506]<=16'd57241;
ROM1[507]<=16'd4730; ROM2[507]<=16'd0; ROM3[507]<=16'd23799; ROM4[507]<=16'd57253;
ROM1[508]<=16'd4764; ROM2[508]<=16'd0; ROM3[508]<=16'd23790; ROM4[508]<=16'd57255;
ROM1[509]<=16'd4778; ROM2[509]<=16'd0; ROM3[509]<=16'd23795; ROM4[509]<=16'd57264;
ROM1[510]<=16'd4771; ROM2[510]<=16'd0; ROM3[510]<=16'd23810; ROM4[510]<=16'd57272;
ROM1[511]<=16'd4748; ROM2[511]<=16'd0; ROM3[511]<=16'd23816; ROM4[511]<=16'd57270;
ROM1[512]<=16'd4726; ROM2[512]<=16'd0; ROM3[512]<=16'd23817; ROM4[512]<=16'd57263;
ROM1[513]<=16'd4707; ROM2[513]<=16'd0; ROM3[513]<=16'd23816; ROM4[513]<=16'd57254;
ROM1[514]<=16'd4719; ROM2[514]<=16'd0; ROM3[514]<=16'd23831; ROM4[514]<=16'd57271;
ROM1[515]<=16'd4731; ROM2[515]<=16'd0; ROM3[515]<=16'd23826; ROM4[515]<=16'd57268;
ROM1[516]<=16'd4742; ROM2[516]<=16'd0; ROM3[516]<=16'd23798; ROM4[516]<=16'd57251;
ROM1[517]<=16'd4753; ROM2[517]<=16'd0; ROM3[517]<=16'd23787; ROM4[517]<=16'd57249;
ROM1[518]<=16'd4738; ROM2[518]<=16'd0; ROM3[518]<=16'd23781; ROM4[518]<=16'd57241;
ROM1[519]<=16'd4721; ROM2[519]<=16'd0; ROM3[519]<=16'd23791; ROM4[519]<=16'd57241;
ROM1[520]<=16'd4715; ROM2[520]<=16'd0; ROM3[520]<=16'd23808; ROM4[520]<=16'd57251;
ROM1[521]<=16'd4705; ROM2[521]<=16'd0; ROM3[521]<=16'd23817; ROM4[521]<=16'd57251;
ROM1[522]<=16'd4708; ROM2[522]<=16'd0; ROM3[522]<=16'd23827; ROM4[522]<=16'd57265;
ROM1[523]<=16'd4728; ROM2[523]<=16'd0; ROM3[523]<=16'd23828; ROM4[523]<=16'd57275;
ROM1[524]<=16'd4744; ROM2[524]<=16'd0; ROM3[524]<=16'd23810; ROM4[524]<=16'd57262;
ROM1[525]<=16'd4771; ROM2[525]<=16'd0; ROM3[525]<=16'd23806; ROM4[525]<=16'd57272;
ROM1[526]<=16'd4755; ROM2[526]<=16'd0; ROM3[526]<=16'd23795; ROM4[526]<=16'd57257;
ROM1[527]<=16'd4738; ROM2[527]<=16'd0; ROM3[527]<=16'd23795; ROM4[527]<=16'd57251;
ROM1[528]<=16'd4752; ROM2[528]<=16'd0; ROM3[528]<=16'd23830; ROM4[528]<=16'd57283;
ROM1[529]<=16'd4736; ROM2[529]<=16'd0; ROM3[529]<=16'd23834; ROM4[529]<=16'd57279;
ROM1[530]<=16'd4710; ROM2[530]<=16'd0; ROM3[530]<=16'd23827; ROM4[530]<=16'd57263;
ROM1[531]<=16'd4717; ROM2[531]<=16'd0; ROM3[531]<=16'd23826; ROM4[531]<=16'd57266;
ROM1[532]<=16'd4735; ROM2[532]<=16'd0; ROM3[532]<=16'd23811; ROM4[532]<=16'd57262;
ROM1[533]<=16'd4772; ROM2[533]<=16'd0; ROM3[533]<=16'd23801; ROM4[533]<=16'd57267;
ROM1[534]<=16'd4783; ROM2[534]<=16'd0; ROM3[534]<=16'd23803; ROM4[534]<=16'd57273;
ROM1[535]<=16'd4761; ROM2[535]<=16'd0; ROM3[535]<=16'd23801; ROM4[535]<=16'd57268;
ROM1[536]<=16'd4731; ROM2[536]<=16'd0; ROM3[536]<=16'd23796; ROM4[536]<=16'd57252;
ROM1[537]<=16'd4707; ROM2[537]<=16'd0; ROM3[537]<=16'd23793; ROM4[537]<=16'd57238;
ROM1[538]<=16'd4695; ROM2[538]<=16'd0; ROM3[538]<=16'd23800; ROM4[538]<=16'd57241;
ROM1[539]<=16'd4692; ROM2[539]<=16'd0; ROM3[539]<=16'd23803; ROM4[539]<=16'd57245;
ROM1[540]<=16'd4710; ROM2[540]<=16'd0; ROM3[540]<=16'd23795; ROM4[540]<=16'd57249;
ROM1[541]<=16'd4750; ROM2[541]<=16'd0; ROM3[541]<=16'd23781; ROM4[541]<=16'd57254;
ROM1[542]<=16'd4769; ROM2[542]<=16'd0; ROM3[542]<=16'd23771; ROM4[542]<=16'd57252;
ROM1[543]<=16'd4755; ROM2[543]<=16'd0; ROM3[543]<=16'd23771; ROM4[543]<=16'd57247;
ROM1[544]<=16'd4735; ROM2[544]<=16'd0; ROM3[544]<=16'd23778; ROM4[544]<=16'd57245;
ROM1[545]<=16'd4713; ROM2[545]<=16'd0; ROM3[545]<=16'd23785; ROM4[545]<=16'd57241;
ROM1[546]<=16'd4702; ROM2[546]<=16'd0; ROM3[546]<=16'd23800; ROM4[546]<=16'd57250;
ROM1[547]<=16'd4703; ROM2[547]<=16'd0; ROM3[547]<=16'd23813; ROM4[547]<=16'd57261;
ROM1[548]<=16'd4712; ROM2[548]<=16'd0; ROM3[548]<=16'd23813; ROM4[548]<=16'd57257;
ROM1[549]<=16'd4740; ROM2[549]<=16'd0; ROM3[549]<=16'd23803; ROM4[549]<=16'd57256;
ROM1[550]<=16'd4765; ROM2[550]<=16'd0; ROM3[550]<=16'd23796; ROM4[550]<=16'd57257;
ROM1[551]<=16'd4763; ROM2[551]<=16'd0; ROM3[551]<=16'd23801; ROM4[551]<=16'd57258;
ROM1[552]<=16'd4747; ROM2[552]<=16'd0; ROM3[552]<=16'd23807; ROM4[552]<=16'd57263;
ROM1[553]<=16'd4717; ROM2[553]<=16'd0; ROM3[553]<=16'd23808; ROM4[553]<=16'd57254;
ROM1[554]<=16'd4699; ROM2[554]<=16'd0; ROM3[554]<=16'd23814; ROM4[554]<=16'd57248;
ROM1[555]<=16'd4689; ROM2[555]<=16'd0; ROM3[555]<=16'd23819; ROM4[555]<=16'd57246;
ROM1[556]<=16'd4700; ROM2[556]<=16'd0; ROM3[556]<=16'd23819; ROM4[556]<=16'd57245;
ROM1[557]<=16'd4733; ROM2[557]<=16'd0; ROM3[557]<=16'd23815; ROM4[557]<=16'd57252;
ROM1[558]<=16'd4759; ROM2[558]<=16'd0; ROM3[558]<=16'd23801; ROM4[558]<=16'd57250;
ROM1[559]<=16'd4757; ROM2[559]<=16'd0; ROM3[559]<=16'd23796; ROM4[559]<=16'd57248;
ROM1[560]<=16'd4743; ROM2[560]<=16'd0; ROM3[560]<=16'd23806; ROM4[560]<=16'd57251;
ROM1[561]<=16'd4728; ROM2[561]<=16'd0; ROM3[561]<=16'd23813; ROM4[561]<=16'd57248;
ROM1[562]<=16'd4714; ROM2[562]<=16'd0; ROM3[562]<=16'd23811; ROM4[562]<=16'd57241;
ROM1[563]<=16'd4698; ROM2[563]<=16'd0; ROM3[563]<=16'd23811; ROM4[563]<=16'd57240;
ROM1[564]<=16'd4699; ROM2[564]<=16'd0; ROM3[564]<=16'd23817; ROM4[564]<=16'd57244;
ROM1[565]<=16'd4716; ROM2[565]<=16'd0; ROM3[565]<=16'd23815; ROM4[565]<=16'd57250;
ROM1[566]<=16'd4746; ROM2[566]<=16'd0; ROM3[566]<=16'd23801; ROM4[566]<=16'd57248;
ROM1[567]<=16'd4767; ROM2[567]<=16'd0; ROM3[567]<=16'd23802; ROM4[567]<=16'd57254;
ROM1[568]<=16'd4761; ROM2[568]<=16'd0; ROM3[568]<=16'd23806; ROM4[568]<=16'd57258;
ROM1[569]<=16'd4748; ROM2[569]<=16'd0; ROM3[569]<=16'd23816; ROM4[569]<=16'd57263;
ROM1[570]<=16'd4729; ROM2[570]<=16'd0; ROM3[570]<=16'd23823; ROM4[570]<=16'd57264;
ROM1[571]<=16'd4712; ROM2[571]<=16'd0; ROM3[571]<=16'd23828; ROM4[571]<=16'd57264;
ROM1[572]<=16'd4699; ROM2[572]<=16'd0; ROM3[572]<=16'd23827; ROM4[572]<=16'd57261;
ROM1[573]<=16'd4712; ROM2[573]<=16'd0; ROM3[573]<=16'd23828; ROM4[573]<=16'd57261;
ROM1[574]<=16'd4756; ROM2[574]<=16'd0; ROM3[574]<=16'd23831; ROM4[574]<=16'd57272;
ROM1[575]<=16'd4785; ROM2[575]<=16'd0; ROM3[575]<=16'd23823; ROM4[575]<=16'd57274;
ROM1[576]<=16'd4788; ROM2[576]<=16'd0; ROM3[576]<=16'd23828; ROM4[576]<=16'd57278;
ROM1[577]<=16'd4772; ROM2[577]<=16'd0; ROM3[577]<=16'd23835; ROM4[577]<=16'd57283;
ROM1[578]<=16'd4766; ROM2[578]<=16'd0; ROM3[578]<=16'd23857; ROM4[578]<=16'd57298;
ROM1[579]<=16'd4766; ROM2[579]<=16'd0; ROM3[579]<=16'd23875; ROM4[579]<=16'd57310;
ROM1[580]<=16'd4738; ROM2[580]<=16'd0; ROM3[580]<=16'd23858; ROM4[580]<=16'd57292;
ROM1[581]<=16'd4714; ROM2[581]<=16'd0; ROM3[581]<=16'd23829; ROM4[581]<=16'd57264;
ROM1[582]<=16'd4728; ROM2[582]<=16'd0; ROM3[582]<=16'd23813; ROM4[582]<=16'd57255;
ROM1[583]<=16'd4755; ROM2[583]<=16'd0; ROM3[583]<=16'd23797; ROM4[583]<=16'd57253;
ROM1[584]<=16'd4773; ROM2[584]<=16'd0; ROM3[584]<=16'd23802; ROM4[584]<=16'd57259;
ROM1[585]<=16'd4780; ROM2[585]<=16'd0; ROM3[585]<=16'd23823; ROM4[585]<=16'd57276;
ROM1[586]<=16'd4770; ROM2[586]<=16'd0; ROM3[586]<=16'd23836; ROM4[586]<=16'd57282;
ROM1[587]<=16'd4751; ROM2[587]<=16'd0; ROM3[587]<=16'd23836; ROM4[587]<=16'd57272;
ROM1[588]<=16'd4723; ROM2[588]<=16'd0; ROM3[588]<=16'd23829; ROM4[588]<=16'd57264;
ROM1[589]<=16'd4719; ROM2[589]<=16'd0; ROM3[589]<=16'd23826; ROM4[589]<=16'd57261;
ROM1[590]<=16'd4721; ROM2[590]<=16'd0; ROM3[590]<=16'd23804; ROM4[590]<=16'd57247;
ROM1[591]<=16'd4747; ROM2[591]<=16'd0; ROM3[591]<=16'd23788; ROM4[591]<=16'd57244;
ROM1[592]<=16'd4762; ROM2[592]<=16'd0; ROM3[592]<=16'd23784; ROM4[592]<=16'd57248;
ROM1[593]<=16'd4751; ROM2[593]<=16'd0; ROM3[593]<=16'd23786; ROM4[593]<=16'd57248;
ROM1[594]<=16'd4740; ROM2[594]<=16'd0; ROM3[594]<=16'd23796; ROM4[594]<=16'd57257;
ROM1[595]<=16'd4731; ROM2[595]<=16'd0; ROM3[595]<=16'd23807; ROM4[595]<=16'd57264;
ROM1[596]<=16'd4719; ROM2[596]<=16'd0; ROM3[596]<=16'd23817; ROM4[596]<=16'd57263;
ROM1[597]<=16'd4708; ROM2[597]<=16'd0; ROM3[597]<=16'd23817; ROM4[597]<=16'd57259;
ROM1[598]<=16'd4718; ROM2[598]<=16'd0; ROM3[598]<=16'd23810; ROM4[598]<=16'd57258;
ROM1[599]<=16'd4741; ROM2[599]<=16'd0; ROM3[599]<=16'd23793; ROM4[599]<=16'd57253;
ROM1[600]<=16'd4767; ROM2[600]<=16'd0; ROM3[600]<=16'd23783; ROM4[600]<=16'd57252;
ROM1[601]<=16'd4759; ROM2[601]<=16'd0; ROM3[601]<=16'd23782; ROM4[601]<=16'd57250;
ROM1[602]<=16'd4733; ROM2[602]<=16'd0; ROM3[602]<=16'd23779; ROM4[602]<=16'd57237;
ROM1[603]<=16'd4718; ROM2[603]<=16'd0; ROM3[603]<=16'd23790; ROM4[603]<=16'd57236;
ROM1[604]<=16'd4711; ROM2[604]<=16'd0; ROM3[604]<=16'd23799; ROM4[604]<=16'd57242;
ROM1[605]<=16'd4702; ROM2[605]<=16'd0; ROM3[605]<=16'd23804; ROM4[605]<=16'd57244;
ROM1[606]<=16'd4713; ROM2[606]<=16'd0; ROM3[606]<=16'd23810; ROM4[606]<=16'd57249;
ROM1[607]<=16'd4746; ROM2[607]<=16'd0; ROM3[607]<=16'd23804; ROM4[607]<=16'd57256;
ROM1[608]<=16'd4786; ROM2[608]<=16'd0; ROM3[608]<=16'd23799; ROM4[608]<=16'd57264;
ROM1[609]<=16'd4796; ROM2[609]<=16'd0; ROM3[609]<=16'd23799; ROM4[609]<=16'd57266;
ROM1[610]<=16'd4761; ROM2[610]<=16'd0; ROM3[610]<=16'd23783; ROM4[610]<=16'd57251;
ROM1[611]<=16'd4729; ROM2[611]<=16'd0; ROM3[611]<=16'd23782; ROM4[611]<=16'd57240;
ROM1[612]<=16'd4713; ROM2[612]<=16'd0; ROM3[612]<=16'd23785; ROM4[612]<=16'd57239;
ROM1[613]<=16'd4699; ROM2[613]<=16'd0; ROM3[613]<=16'd23794; ROM4[613]<=16'd57245;
ROM1[614]<=16'd4710; ROM2[614]<=16'd0; ROM3[614]<=16'd23808; ROM4[614]<=16'd57257;
ROM1[615]<=16'd4734; ROM2[615]<=16'd0; ROM3[615]<=16'd23799; ROM4[615]<=16'd57257;
ROM1[616]<=16'd4761; ROM2[616]<=16'd0; ROM3[616]<=16'd23779; ROM4[616]<=16'd57251;
ROM1[617]<=16'd4784; ROM2[617]<=16'd0; ROM3[617]<=16'd23782; ROM4[617]<=16'd57259;
ROM1[618]<=16'd4779; ROM2[618]<=16'd0; ROM3[618]<=16'd23795; ROM4[618]<=16'd57267;
ROM1[619]<=16'd4761; ROM2[619]<=16'd0; ROM3[619]<=16'd23809; ROM4[619]<=16'd57272;
ROM1[620]<=16'd4759; ROM2[620]<=16'd0; ROM3[620]<=16'd23830; ROM4[620]<=16'd57282;
ROM1[621]<=16'd4729; ROM2[621]<=16'd0; ROM3[621]<=16'd23826; ROM4[621]<=16'd57268;
ROM1[622]<=16'd4702; ROM2[622]<=16'd0; ROM3[622]<=16'd23812; ROM4[622]<=16'd57255;
ROM1[623]<=16'd4714; ROM2[623]<=16'd0; ROM3[623]<=16'd23809; ROM4[623]<=16'd57254;
ROM1[624]<=16'd4741; ROM2[624]<=16'd0; ROM3[624]<=16'd23797; ROM4[624]<=16'd57251;
ROM1[625]<=16'd4772; ROM2[625]<=16'd0; ROM3[625]<=16'd23790; ROM4[625]<=16'd57258;
ROM1[626]<=16'd4781; ROM2[626]<=16'd0; ROM3[626]<=16'd23799; ROM4[626]<=16'd57269;
ROM1[627]<=16'd4750; ROM2[627]<=16'd0; ROM3[627]<=16'd23796; ROM4[627]<=16'd57258;
ROM1[628]<=16'd4719; ROM2[628]<=16'd0; ROM3[628]<=16'd23796; ROM4[628]<=16'd57250;
ROM1[629]<=16'd4712; ROM2[629]<=16'd0; ROM3[629]<=16'd23807; ROM4[629]<=16'd57256;
ROM1[630]<=16'd4707; ROM2[630]<=16'd0; ROM3[630]<=16'd23813; ROM4[630]<=16'd57255;
ROM1[631]<=16'd4725; ROM2[631]<=16'd0; ROM3[631]<=16'd23825; ROM4[631]<=16'd57269;
ROM1[632]<=16'd4762; ROM2[632]<=16'd0; ROM3[632]<=16'd23830; ROM4[632]<=16'd57281;
ROM1[633]<=16'd4789; ROM2[633]<=16'd0; ROM3[633]<=16'd23813; ROM4[633]<=16'd57279;
ROM1[634]<=16'd4793; ROM2[634]<=16'd0; ROM3[634]<=16'd23808; ROM4[634]<=16'd57284;
ROM1[635]<=16'd4775; ROM2[635]<=16'd0; ROM3[635]<=16'd23810; ROM4[635]<=16'd57284;
ROM1[636]<=16'd4740; ROM2[636]<=16'd0; ROM3[636]<=16'd23806; ROM4[636]<=16'd57268;
ROM1[637]<=16'd4718; ROM2[637]<=16'd0; ROM3[637]<=16'd23808; ROM4[637]<=16'd57260;
ROM1[638]<=16'd4707; ROM2[638]<=16'd0; ROM3[638]<=16'd23818; ROM4[638]<=16'd57261;
ROM1[639]<=16'd4712; ROM2[639]<=16'd0; ROM3[639]<=16'd23821; ROM4[639]<=16'd57265;
ROM1[640]<=16'd4735; ROM2[640]<=16'd0; ROM3[640]<=16'd23819; ROM4[640]<=16'd57273;
ROM1[641]<=16'd4781; ROM2[641]<=16'd0; ROM3[641]<=16'd23818; ROM4[641]<=16'd57290;
ROM1[642]<=16'd4796; ROM2[642]<=16'd0; ROM3[642]<=16'd23807; ROM4[642]<=16'd57286;
ROM1[643]<=16'd4769; ROM2[643]<=16'd0; ROM3[643]<=16'd23788; ROM4[643]<=16'd57264;
ROM1[644]<=16'd4750; ROM2[644]<=16'd0; ROM3[644]<=16'd23786; ROM4[644]<=16'd57258;
ROM1[645]<=16'd4734; ROM2[645]<=16'd0; ROM3[645]<=16'd23792; ROM4[645]<=16'd57258;
ROM1[646]<=16'd4719; ROM2[646]<=16'd0; ROM3[646]<=16'd23802; ROM4[646]<=16'd57261;
ROM1[647]<=16'd4717; ROM2[647]<=16'd0; ROM3[647]<=16'd23810; ROM4[647]<=16'd57266;
ROM1[648]<=16'd4718; ROM2[648]<=16'd0; ROM3[648]<=16'd23795; ROM4[648]<=16'd57258;
ROM1[649]<=16'd4741; ROM2[649]<=16'd0; ROM3[649]<=16'd23777; ROM4[649]<=16'd57250;
ROM1[650]<=16'd4767; ROM2[650]<=16'd0; ROM3[650]<=16'd23771; ROM4[650]<=16'd57249;
ROM1[651]<=16'd4764; ROM2[651]<=16'd0; ROM3[651]<=16'd23772; ROM4[651]<=16'd57252;
ROM1[652]<=16'd4759; ROM2[652]<=16'd0; ROM3[652]<=16'd23791; ROM4[652]<=16'd57264;
ROM1[653]<=16'd4738; ROM2[653]<=16'd0; ROM3[653]<=16'd23800; ROM4[653]<=16'd57259;
ROM1[654]<=16'd4721; ROM2[654]<=16'd0; ROM3[654]<=16'd23797; ROM4[654]<=16'd57253;
ROM1[655]<=16'd4728; ROM2[655]<=16'd0; ROM3[655]<=16'd23820; ROM4[655]<=16'd57267;
ROM1[656]<=16'd4741; ROM2[656]<=16'd0; ROM3[656]<=16'd23830; ROM4[656]<=16'd57275;
ROM1[657]<=16'd4763; ROM2[657]<=16'd0; ROM3[657]<=16'd23814; ROM4[657]<=16'd57269;
ROM1[658]<=16'd4789; ROM2[658]<=16'd0; ROM3[658]<=16'd23796; ROM4[658]<=16'd57263;
ROM1[659]<=16'd4793; ROM2[659]<=16'd0; ROM3[659]<=16'd23797; ROM4[659]<=16'd57265;
ROM1[660]<=16'd4764; ROM2[660]<=16'd0; ROM3[660]<=16'd23795; ROM4[660]<=16'd57257;
ROM1[661]<=16'd4739; ROM2[661]<=16'd0; ROM3[661]<=16'd23798; ROM4[661]<=16'd57253;
ROM1[662]<=16'd4737; ROM2[662]<=16'd0; ROM3[662]<=16'd23816; ROM4[662]<=16'd57268;
ROM1[663]<=16'd4729; ROM2[663]<=16'd0; ROM3[663]<=16'd23825; ROM4[663]<=16'd57268;
ROM1[664]<=16'd4722; ROM2[664]<=16'd0; ROM3[664]<=16'd23811; ROM4[664]<=16'd57257;
ROM1[665]<=16'd4731; ROM2[665]<=16'd0; ROM3[665]<=16'd23794; ROM4[665]<=16'd57251;
ROM1[666]<=16'd4756; ROM2[666]<=16'd0; ROM3[666]<=16'd23771; ROM4[666]<=16'd57239;
ROM1[667]<=16'd4761; ROM2[667]<=16'd0; ROM3[667]<=16'd23753; ROM4[667]<=16'd57231;
ROM1[668]<=16'd4749; ROM2[668]<=16'd0; ROM3[668]<=16'd23762; ROM4[668]<=16'd57236;
ROM1[669]<=16'd4734; ROM2[669]<=16'd0; ROM3[669]<=16'd23779; ROM4[669]<=16'd57245;
ROM1[670]<=16'd4723; ROM2[670]<=16'd0; ROM3[670]<=16'd23791; ROM4[670]<=16'd57252;
ROM1[671]<=16'd4707; ROM2[671]<=16'd0; ROM3[671]<=16'd23793; ROM4[671]<=16'd57246;
ROM1[672]<=16'd4705; ROM2[672]<=16'd0; ROM3[672]<=16'd23793; ROM4[672]<=16'd57247;
ROM1[673]<=16'd4725; ROM2[673]<=16'd0; ROM3[673]<=16'd23794; ROM4[673]<=16'd57250;
ROM1[674]<=16'd4738; ROM2[674]<=16'd0; ROM3[674]<=16'd23775; ROM4[674]<=16'd57234;
ROM1[675]<=16'd4749; ROM2[675]<=16'd0; ROM3[675]<=16'd23761; ROM4[675]<=16'd57228;
ROM1[676]<=16'd4751; ROM2[676]<=16'd0; ROM3[676]<=16'd23766; ROM4[676]<=16'd57231;
ROM1[677]<=16'd4734; ROM2[677]<=16'd0; ROM3[677]<=16'd23769; ROM4[677]<=16'd57227;
ROM1[678]<=16'd4711; ROM2[678]<=16'd0; ROM3[678]<=16'd23767; ROM4[678]<=16'd57220;
ROM1[679]<=16'd4690; ROM2[679]<=16'd0; ROM3[679]<=16'd23769; ROM4[679]<=16'd57216;
ROM1[680]<=16'd4676; ROM2[680]<=16'd0; ROM3[680]<=16'd23775; ROM4[680]<=16'd57213;
ROM1[681]<=16'd4680; ROM2[681]<=16'd0; ROM3[681]<=16'd23774; ROM4[681]<=16'd57209;
ROM1[682]<=16'd4716; ROM2[682]<=16'd0; ROM3[682]<=16'd23775; ROM4[682]<=16'd57219;
ROM1[683]<=16'd4763; ROM2[683]<=16'd0; ROM3[683]<=16'd23773; ROM4[683]<=16'd57235;
ROM1[684]<=16'd4772; ROM2[684]<=16'd0; ROM3[684]<=16'd23778; ROM4[684]<=16'd57241;
ROM1[685]<=16'd4752; ROM2[685]<=16'd0; ROM3[685]<=16'd23783; ROM4[685]<=16'd57243;
ROM1[686]<=16'd4755; ROM2[686]<=16'd0; ROM3[686]<=16'd23814; ROM4[686]<=16'd57269;
ROM1[687]<=16'd4767; ROM2[687]<=16'd0; ROM3[687]<=16'd23846; ROM4[687]<=16'd57291;
ROM1[688]<=16'd4727; ROM2[688]<=16'd0; ROM3[688]<=16'd23821; ROM4[688]<=16'd57266;
ROM1[689]<=16'd4704; ROM2[689]<=16'd0; ROM3[689]<=16'd23799; ROM4[689]<=16'd57246;
ROM1[690]<=16'd4718; ROM2[690]<=16'd0; ROM3[690]<=16'd23791; ROM4[690]<=16'd57243;
ROM1[691]<=16'd4738; ROM2[691]<=16'd0; ROM3[691]<=16'd23774; ROM4[691]<=16'd57236;
ROM1[692]<=16'd4760; ROM2[692]<=16'd0; ROM3[692]<=16'd23780; ROM4[692]<=16'd57245;
ROM1[693]<=16'd4767; ROM2[693]<=16'd0; ROM3[693]<=16'd23802; ROM4[693]<=16'd57266;
ROM1[694]<=16'd4749; ROM2[694]<=16'd0; ROM3[694]<=16'd23812; ROM4[694]<=16'd57270;
ROM1[695]<=16'd4741; ROM2[695]<=16'd0; ROM3[695]<=16'd23824; ROM4[695]<=16'd57276;
ROM1[696]<=16'd4740; ROM2[696]<=16'd0; ROM3[696]<=16'd23839; ROM4[696]<=16'd57292;
ROM1[697]<=16'd4735; ROM2[697]<=16'd0; ROM3[697]<=16'd23844; ROM4[697]<=16'd57294;
ROM1[698]<=16'd4743; ROM2[698]<=16'd0; ROM3[698]<=16'd23839; ROM4[698]<=16'd57292;
ROM1[699]<=16'd4766; ROM2[699]<=16'd0; ROM3[699]<=16'd23821; ROM4[699]<=16'd57284;
ROM1[700]<=16'd4810; ROM2[700]<=16'd0; ROM3[700]<=16'd23829; ROM4[700]<=16'd57299;
ROM1[701]<=16'd4814; ROM2[701]<=16'd0; ROM3[701]<=16'd23833; ROM4[701]<=16'd57307;
ROM1[702]<=16'd4780; ROM2[702]<=16'd0; ROM3[702]<=16'd23815; ROM4[702]<=16'd57286;
ROM1[703]<=16'd4756; ROM2[703]<=16'd0; ROM3[703]<=16'd23811; ROM4[703]<=16'd57275;
ROM1[704]<=16'd4744; ROM2[704]<=16'd0; ROM3[704]<=16'd23817; ROM4[704]<=16'd57275;
ROM1[705]<=16'd4731; ROM2[705]<=16'd0; ROM3[705]<=16'd23826; ROM4[705]<=16'd57272;
ROM1[706]<=16'd4734; ROM2[706]<=16'd0; ROM3[706]<=16'd23819; ROM4[706]<=16'd57266;
ROM1[707]<=16'd4757; ROM2[707]<=16'd0; ROM3[707]<=16'd23807; ROM4[707]<=16'd57270;
ROM1[708]<=16'd4785; ROM2[708]<=16'd0; ROM3[708]<=16'd23792; ROM4[708]<=16'd57269;
ROM1[709]<=16'd4795; ROM2[709]<=16'd0; ROM3[709]<=16'd23793; ROM4[709]<=16'd57271;
ROM1[710]<=16'd4791; ROM2[710]<=16'd0; ROM3[710]<=16'd23809; ROM4[710]<=16'd57284;
ROM1[711]<=16'd4780; ROM2[711]<=16'd0; ROM3[711]<=16'd23821; ROM4[711]<=16'd57293;
ROM1[712]<=16'd4763; ROM2[712]<=16'd0; ROM3[712]<=16'd23823; ROM4[712]<=16'd57291;
ROM1[713]<=16'd4742; ROM2[713]<=16'd0; ROM3[713]<=16'd23823; ROM4[713]<=16'd57282;
ROM1[714]<=16'd4737; ROM2[714]<=16'd0; ROM3[714]<=16'd23820; ROM4[714]<=16'd57279;
ROM1[715]<=16'd4745; ROM2[715]<=16'd0; ROM3[715]<=16'd23807; ROM4[715]<=16'd57271;
ROM1[716]<=16'd4768; ROM2[716]<=16'd0; ROM3[716]<=16'd23783; ROM4[716]<=16'd57262;
ROM1[717]<=16'd4779; ROM2[717]<=16'd0; ROM3[717]<=16'd23769; ROM4[717]<=16'd57258;
ROM1[718]<=16'd4766; ROM2[718]<=16'd0; ROM3[718]<=16'd23768; ROM4[718]<=16'd57255;
ROM1[719]<=16'd4748; ROM2[719]<=16'd0; ROM3[719]<=16'd23769; ROM4[719]<=16'd57248;
ROM1[720]<=16'd4728; ROM2[720]<=16'd0; ROM3[720]<=16'd23772; ROM4[720]<=16'd57241;
ROM1[721]<=16'd4708; ROM2[721]<=16'd0; ROM3[721]<=16'd23782; ROM4[721]<=16'd57239;
ROM1[722]<=16'd4699; ROM2[722]<=16'd0; ROM3[722]<=16'd23785; ROM4[722]<=16'd57240;
ROM1[723]<=16'd4710; ROM2[723]<=16'd0; ROM3[723]<=16'd23783; ROM4[723]<=16'd57240;
ROM1[724]<=16'd4741; ROM2[724]<=16'd0; ROM3[724]<=16'd23778; ROM4[724]<=16'd57242;
ROM1[725]<=16'd4777; ROM2[725]<=16'd0; ROM3[725]<=16'd23772; ROM4[725]<=16'd57252;
ROM1[726]<=16'd4779; ROM2[726]<=16'd0; ROM3[726]<=16'd23775; ROM4[726]<=16'd57257;
ROM1[727]<=16'd4757; ROM2[727]<=16'd0; ROM3[727]<=16'd23778; ROM4[727]<=16'd57253;
ROM1[728]<=16'd4736; ROM2[728]<=16'd0; ROM3[728]<=16'd23789; ROM4[728]<=16'd57251;
ROM1[729]<=16'd4730; ROM2[729]<=16'd0; ROM3[729]<=16'd23808; ROM4[729]<=16'd57263;
ROM1[730]<=16'd4726; ROM2[730]<=16'd0; ROM3[730]<=16'd23829; ROM4[730]<=16'd57274;
ROM1[731]<=16'd4728; ROM2[731]<=16'd0; ROM3[731]<=16'd23822; ROM4[731]<=16'd57268;
ROM1[732]<=16'd4747; ROM2[732]<=16'd0; ROM3[732]<=16'd23805; ROM4[732]<=16'd57258;
ROM1[733]<=16'd4767; ROM2[733]<=16'd0; ROM3[733]<=16'd23784; ROM4[733]<=16'd57249;
ROM1[734]<=16'd4768; ROM2[734]<=16'd0; ROM3[734]<=16'd23780; ROM4[734]<=16'd57249;
ROM1[735]<=16'd4765; ROM2[735]<=16'd0; ROM3[735]<=16'd23802; ROM4[735]<=16'd57262;
ROM1[736]<=16'd4773; ROM2[736]<=16'd0; ROM3[736]<=16'd23837; ROM4[736]<=16'd57289;
ROM1[737]<=16'd4787; ROM2[737]<=16'd0; ROM3[737]<=16'd23865; ROM4[737]<=16'd57310;
ROM1[738]<=16'd4767; ROM2[738]<=16'd0; ROM3[738]<=16'd23859; ROM4[738]<=16'd57299;
ROM1[739]<=16'd4739; ROM2[739]<=16'd0; ROM3[739]<=16'd23839; ROM4[739]<=16'd57275;
ROM1[740]<=16'd4739; ROM2[740]<=16'd0; ROM3[740]<=16'd23816; ROM4[740]<=16'd57258;
ROM1[741]<=16'd4765; ROM2[741]<=16'd0; ROM3[741]<=16'd23800; ROM4[741]<=16'd57256;
ROM1[742]<=16'd4800; ROM2[742]<=16'd0; ROM3[742]<=16'd23812; ROM4[742]<=16'd57276;
ROM1[743]<=16'd4805; ROM2[743]<=16'd0; ROM3[743]<=16'd23831; ROM4[743]<=16'd57290;
ROM1[744]<=16'd4771; ROM2[744]<=16'd0; ROM3[744]<=16'd23828; ROM4[744]<=16'd57278;
ROM1[745]<=16'd4751; ROM2[745]<=16'd0; ROM3[745]<=16'd23830; ROM4[745]<=16'd57274;
ROM1[746]<=16'd4732; ROM2[746]<=16'd0; ROM3[746]<=16'd23833; ROM4[746]<=16'd57274;
ROM1[747]<=16'd4731; ROM2[747]<=16'd0; ROM3[747]<=16'd23837; ROM4[747]<=16'd57283;
ROM1[748]<=16'd4768; ROM2[748]<=16'd0; ROM3[748]<=16'd23853; ROM4[748]<=16'd57304;
ROM1[749]<=16'd4792; ROM2[749]<=16'd0; ROM3[749]<=16'd23837; ROM4[749]<=16'd57295;
ROM1[750]<=16'd4807; ROM2[750]<=16'd0; ROM3[750]<=16'd23818; ROM4[750]<=16'd57283;
ROM1[751]<=16'd4816; ROM2[751]<=16'd0; ROM3[751]<=16'd23835; ROM4[751]<=16'd57301;
ROM1[752]<=16'd4796; ROM2[752]<=16'd0; ROM3[752]<=16'd23838; ROM4[752]<=16'd57301;
ROM1[753]<=16'd4777; ROM2[753]<=16'd0; ROM3[753]<=16'd23839; ROM4[753]<=16'd57295;
ROM1[754]<=16'd4767; ROM2[754]<=16'd0; ROM3[754]<=16'd23847; ROM4[754]<=16'd57295;
ROM1[755]<=16'd4749; ROM2[755]<=16'd0; ROM3[755]<=16'd23843; ROM4[755]<=16'd57286;
ROM1[756]<=16'd4754; ROM2[756]<=16'd0; ROM3[756]<=16'd23839; ROM4[756]<=16'd57288;
ROM1[757]<=16'd4781; ROM2[757]<=16'd0; ROM3[757]<=16'd23836; ROM4[757]<=16'd57294;
ROM1[758]<=16'd4813; ROM2[758]<=16'd0; ROM3[758]<=16'd23832; ROM4[758]<=16'd57298;
ROM1[759]<=16'd4820; ROM2[759]<=16'd0; ROM3[759]<=16'd23835; ROM4[759]<=16'd57303;
ROM1[760]<=16'd4797; ROM2[760]<=16'd0; ROM3[760]<=16'd23834; ROM4[760]<=16'd57293;
ROM1[761]<=16'd4775; ROM2[761]<=16'd0; ROM3[761]<=16'd23837; ROM4[761]<=16'd57292;
ROM1[762]<=16'd4770; ROM2[762]<=16'd0; ROM3[762]<=16'd23850; ROM4[762]<=16'd57302;
ROM1[763]<=16'd4744; ROM2[763]<=16'd0; ROM3[763]<=16'd23840; ROM4[763]<=16'd57283;
ROM1[764]<=16'd4733; ROM2[764]<=16'd0; ROM3[764]<=16'd23828; ROM4[764]<=16'd57274;
ROM1[765]<=16'd4748; ROM2[765]<=16'd0; ROM3[765]<=16'd23814; ROM4[765]<=16'd57270;
ROM1[766]<=16'd4770; ROM2[766]<=16'd0; ROM3[766]<=16'd23791; ROM4[766]<=16'd57254;
ROM1[767]<=16'd4778; ROM2[767]<=16'd0; ROM3[767]<=16'd23775; ROM4[767]<=16'd57247;
ROM1[768]<=16'd4765; ROM2[768]<=16'd0; ROM3[768]<=16'd23781; ROM4[768]<=16'd57247;
ROM1[769]<=16'd4755; ROM2[769]<=16'd0; ROM3[769]<=16'd23797; ROM4[769]<=16'd57252;
ROM1[770]<=16'd4739; ROM2[770]<=16'd0; ROM3[770]<=16'd23800; ROM4[770]<=16'd57249;
ROM1[771]<=16'd4721; ROM2[771]<=16'd0; ROM3[771]<=16'd23807; ROM4[771]<=16'd57248;
ROM1[772]<=16'd4732; ROM2[772]<=16'd0; ROM3[772]<=16'd23829; ROM4[772]<=16'd57266;
ROM1[773]<=16'd4765; ROM2[773]<=16'd0; ROM3[773]<=16'd23850; ROM4[773]<=16'd57288;
ROM1[774]<=16'd4793; ROM2[774]<=16'd0; ROM3[774]<=16'd23842; ROM4[774]<=16'd57290;
ROM1[775]<=16'd4806; ROM2[775]<=16'd0; ROM3[775]<=16'd23820; ROM4[775]<=16'd57283;
ROM1[776]<=16'd4788; ROM2[776]<=16'd0; ROM3[776]<=16'd23811; ROM4[776]<=16'd57274;
ROM1[777]<=16'd4753; ROM2[777]<=16'd0; ROM3[777]<=16'd23803; ROM4[777]<=16'd57259;
ROM1[778]<=16'd4729; ROM2[778]<=16'd0; ROM3[778]<=16'd23800; ROM4[778]<=16'd57251;
ROM1[779]<=16'd4726; ROM2[779]<=16'd0; ROM3[779]<=16'd23820; ROM4[779]<=16'd57265;
ROM1[780]<=16'd4721; ROM2[780]<=16'd0; ROM3[780]<=16'd23832; ROM4[780]<=16'd57273;
ROM1[781]<=16'd4721; ROM2[781]<=16'd0; ROM3[781]<=16'd23822; ROM4[781]<=16'd57265;
ROM1[782]<=16'd4745; ROM2[782]<=16'd0; ROM3[782]<=16'd23813; ROM4[782]<=16'd57265;
ROM1[783]<=16'd4778; ROM2[783]<=16'd0; ROM3[783]<=16'd23800; ROM4[783]<=16'd57263;
ROM1[784]<=16'd4789; ROM2[784]<=16'd0; ROM3[784]<=16'd23803; ROM4[784]<=16'd57271;
ROM1[785]<=16'd4777; ROM2[785]<=16'd0; ROM3[785]<=16'd23815; ROM4[785]<=16'd57277;
ROM1[786]<=16'd4761; ROM2[786]<=16'd0; ROM3[786]<=16'd23823; ROM4[786]<=16'd57282;
ROM1[787]<=16'd4756; ROM2[787]<=16'd0; ROM3[787]<=16'd23838; ROM4[787]<=16'd57291;
ROM1[788]<=16'd4750; ROM2[788]<=16'd0; ROM3[788]<=16'd23846; ROM4[788]<=16'd57293;
ROM1[789]<=16'd4741; ROM2[789]<=16'd0; ROM3[789]<=16'd23833; ROM4[789]<=16'd57279;
ROM1[790]<=16'd4751; ROM2[790]<=16'd0; ROM3[790]<=16'd23817; ROM4[790]<=16'd57271;
ROM1[791]<=16'd4782; ROM2[791]<=16'd0; ROM3[791]<=16'd23802; ROM4[791]<=16'd57271;
ROM1[792]<=16'd4792; ROM2[792]<=16'd0; ROM3[792]<=16'd23784; ROM4[792]<=16'd57260;
ROM1[793]<=16'd4776; ROM2[793]<=16'd0; ROM3[793]<=16'd23786; ROM4[793]<=16'd57263;
ROM1[794]<=16'd4758; ROM2[794]<=16'd0; ROM3[794]<=16'd23799; ROM4[794]<=16'd57267;
ROM1[795]<=16'd4742; ROM2[795]<=16'd0; ROM3[795]<=16'd23805; ROM4[795]<=16'd57262;
ROM1[796]<=16'd4724; ROM2[796]<=16'd0; ROM3[796]<=16'd23812; ROM4[796]<=16'd57264;
ROM1[797]<=16'd4724; ROM2[797]<=16'd0; ROM3[797]<=16'd23820; ROM4[797]<=16'd57268;
ROM1[798]<=16'd4739; ROM2[798]<=16'd0; ROM3[798]<=16'd23819; ROM4[798]<=16'd57265;
ROM1[799]<=16'd4769; ROM2[799]<=16'd0; ROM3[799]<=16'd23810; ROM4[799]<=16'd57267;
ROM1[800]<=16'd4784; ROM2[800]<=16'd0; ROM3[800]<=16'd23794; ROM4[800]<=16'd57260;
ROM1[801]<=16'd4768; ROM2[801]<=16'd0; ROM3[801]<=16'd23784; ROM4[801]<=16'd57248;
ROM1[802]<=16'd4753; ROM2[802]<=16'd0; ROM3[802]<=16'd23793; ROM4[802]<=16'd57250;
ROM1[803]<=16'd4736; ROM2[803]<=16'd0; ROM3[803]<=16'd23799; ROM4[803]<=16'd57250;
ROM1[804]<=16'd4725; ROM2[804]<=16'd0; ROM3[804]<=16'd23811; ROM4[804]<=16'd57258;
ROM1[805]<=16'd4718; ROM2[805]<=16'd0; ROM3[805]<=16'd23822; ROM4[805]<=16'd57265;
ROM1[806]<=16'd4718; ROM2[806]<=16'd0; ROM3[806]<=16'd23814; ROM4[806]<=16'd57264;
ROM1[807]<=16'd4740; ROM2[807]<=16'd0; ROM3[807]<=16'd23810; ROM4[807]<=16'd57265;
ROM1[808]<=16'd4771; ROM2[808]<=16'd0; ROM3[808]<=16'd23795; ROM4[808]<=16'd57262;
ROM1[809]<=16'd4777; ROM2[809]<=16'd0; ROM3[809]<=16'd23793; ROM4[809]<=16'd57265;
ROM1[810]<=16'd4766; ROM2[810]<=16'd0; ROM3[810]<=16'd23807; ROM4[810]<=16'd57272;
ROM1[811]<=16'd4758; ROM2[811]<=16'd0; ROM3[811]<=16'd23820; ROM4[811]<=16'd57281;
ROM1[812]<=16'd4754; ROM2[812]<=16'd0; ROM3[812]<=16'd23829; ROM4[812]<=16'd57292;
ROM1[813]<=16'd4748; ROM2[813]<=16'd0; ROM3[813]<=16'd23841; ROM4[813]<=16'd57300;
ROM1[814]<=16'd4748; ROM2[814]<=16'd0; ROM3[814]<=16'd23843; ROM4[814]<=16'd57299;
ROM1[815]<=16'd4756; ROM2[815]<=16'd0; ROM3[815]<=16'd23830; ROM4[815]<=16'd57291;
ROM1[816]<=16'd4781; ROM2[816]<=16'd0; ROM3[816]<=16'd23815; ROM4[816]<=16'd57282;
ROM1[817]<=16'd4779; ROM2[817]<=16'd0; ROM3[817]<=16'd23792; ROM4[817]<=16'd57271;
ROM1[818]<=16'd4754; ROM2[818]<=16'd0; ROM3[818]<=16'd23784; ROM4[818]<=16'd57258;
ROM1[819]<=16'd4741; ROM2[819]<=16'd0; ROM3[819]<=16'd23793; ROM4[819]<=16'd57259;
ROM1[820]<=16'd4733; ROM2[820]<=16'd0; ROM3[820]<=16'd23809; ROM4[820]<=16'd57265;
ROM1[821]<=16'd4723; ROM2[821]<=16'd0; ROM3[821]<=16'd23827; ROM4[821]<=16'd57271;
ROM1[822]<=16'd4719; ROM2[822]<=16'd0; ROM3[822]<=16'd23832; ROM4[822]<=16'd57278;
ROM1[823]<=16'd4733; ROM2[823]<=16'd0; ROM3[823]<=16'd23827; ROM4[823]<=16'd57279;
ROM1[824]<=16'd4769; ROM2[824]<=16'd0; ROM3[824]<=16'd23826; ROM4[824]<=16'd57287;
ROM1[825]<=16'd4787; ROM2[825]<=16'd0; ROM3[825]<=16'd23816; ROM4[825]<=16'd57283;
ROM1[826]<=16'd4772; ROM2[826]<=16'd0; ROM3[826]<=16'd23811; ROM4[826]<=16'd57274;
ROM1[827]<=16'd4755; ROM2[827]<=16'd0; ROM3[827]<=16'd23822; ROM4[827]<=16'd57277;
ROM1[828]<=16'd4723; ROM2[828]<=16'd0; ROM3[828]<=16'd23820; ROM4[828]<=16'd57265;
ROM1[829]<=16'd4704; ROM2[829]<=16'd0; ROM3[829]<=16'd23820; ROM4[829]<=16'd57258;
ROM1[830]<=16'd4709; ROM2[830]<=16'd0; ROM3[830]<=16'd23836; ROM4[830]<=16'd57270;
ROM1[831]<=16'd4743; ROM2[831]<=16'd0; ROM3[831]<=16'd23860; ROM4[831]<=16'd57295;
ROM1[832]<=16'd4765; ROM2[832]<=16'd0; ROM3[832]<=16'd23843; ROM4[832]<=16'd57293;
ROM1[833]<=16'd4779; ROM2[833]<=16'd0; ROM3[833]<=16'd23814; ROM4[833]<=16'd57277;
ROM1[834]<=16'd4786; ROM2[834]<=16'd0; ROM3[834]<=16'd23814; ROM4[834]<=16'd57276;
ROM1[835]<=16'd4766; ROM2[835]<=16'd0; ROM3[835]<=16'd23815; ROM4[835]<=16'd57276;
ROM1[836]<=16'd4754; ROM2[836]<=16'd0; ROM3[836]<=16'd23832; ROM4[836]<=16'd57284;
ROM1[837]<=16'd4749; ROM2[837]<=16'd0; ROM3[837]<=16'd23838; ROM4[837]<=16'd57288;
ROM1[838]<=16'd4719; ROM2[838]<=16'd0; ROM3[838]<=16'd23825; ROM4[838]<=16'd57275;
ROM1[839]<=16'd4703; ROM2[839]<=16'd0; ROM3[839]<=16'd23811; ROM4[839]<=16'd57261;
ROM1[840]<=16'd4707; ROM2[840]<=16'd0; ROM3[840]<=16'd23786; ROM4[840]<=16'd57246;
ROM1[841]<=16'd4737; ROM2[841]<=16'd0; ROM3[841]<=16'd23773; ROM4[841]<=16'd57245;
ROM1[842]<=16'd4765; ROM2[842]<=16'd0; ROM3[842]<=16'd23785; ROM4[842]<=16'd57260;
ROM1[843]<=16'd4755; ROM2[843]<=16'd0; ROM3[843]<=16'd23791; ROM4[843]<=16'd57261;
ROM1[844]<=16'd4729; ROM2[844]<=16'd0; ROM3[844]<=16'd23792; ROM4[844]<=16'd57256;
ROM1[845]<=16'd4710; ROM2[845]<=16'd0; ROM3[845]<=16'd23798; ROM4[845]<=16'd57252;
ROM1[846]<=16'd4714; ROM2[846]<=16'd0; ROM3[846]<=16'd23820; ROM4[846]<=16'd57272;
ROM1[847]<=16'd4705; ROM2[847]<=16'd0; ROM3[847]<=16'd23821; ROM4[847]<=16'd57270;
ROM1[848]<=16'd4711; ROM2[848]<=16'd0; ROM3[848]<=16'd23808; ROM4[848]<=16'd57258;
ROM1[849]<=16'd4746; ROM2[849]<=16'd0; ROM3[849]<=16'd23801; ROM4[849]<=16'd57265;
ROM1[850]<=16'd4766; ROM2[850]<=16'd0; ROM3[850]<=16'd23790; ROM4[850]<=16'd57266;
ROM1[851]<=16'd4752; ROM2[851]<=16'd0; ROM3[851]<=16'd23780; ROM4[851]<=16'd57257;
ROM1[852]<=16'd4741; ROM2[852]<=16'd0; ROM3[852]<=16'd23791; ROM4[852]<=16'd57261;
ROM1[853]<=16'd4744; ROM2[853]<=16'd0; ROM3[853]<=16'd23818; ROM4[853]<=16'd57276;
ROM1[854]<=16'd4722; ROM2[854]<=16'd0; ROM3[854]<=16'd23819; ROM4[854]<=16'd57272;
ROM1[855]<=16'd4708; ROM2[855]<=16'd0; ROM3[855]<=16'd23830; ROM4[855]<=16'd57273;
ROM1[856]<=16'd4718; ROM2[856]<=16'd0; ROM3[856]<=16'd23843; ROM4[856]<=16'd57283;
ROM1[857]<=16'd4748; ROM2[857]<=16'd0; ROM3[857]<=16'd23841; ROM4[857]<=16'd57291;
ROM1[858]<=16'd4781; ROM2[858]<=16'd0; ROM3[858]<=16'd23833; ROM4[858]<=16'd57293;
ROM1[859]<=16'd4793; ROM2[859]<=16'd0; ROM3[859]<=16'd23837; ROM4[859]<=16'd57298;
ROM1[860]<=16'd4794; ROM2[860]<=16'd0; ROM3[860]<=16'd23861; ROM4[860]<=16'd57313;
ROM1[861]<=16'd4772; ROM2[861]<=16'd0; ROM3[861]<=16'd23872; ROM4[861]<=16'd57314;
ROM1[862]<=16'd4757; ROM2[862]<=16'd0; ROM3[862]<=16'd23874; ROM4[862]<=16'd57311;
ROM1[863]<=16'd4745; ROM2[863]<=16'd0; ROM3[863]<=16'd23879; ROM4[863]<=16'd57315;
ROM1[864]<=16'd4739; ROM2[864]<=16'd0; ROM3[864]<=16'd23872; ROM4[864]<=16'd57315;
ROM1[865]<=16'd4780; ROM2[865]<=16'd0; ROM3[865]<=16'd23879; ROM4[865]<=16'd57337;
ROM1[866]<=16'd4821; ROM2[866]<=16'd0; ROM3[866]<=16'd23872; ROM4[866]<=16'd57339;
ROM1[867]<=16'd4812; ROM2[867]<=16'd0; ROM3[867]<=16'd23845; ROM4[867]<=16'd57319;
ROM1[868]<=16'd4788; ROM2[868]<=16'd0; ROM3[868]<=16'd23840; ROM4[868]<=16'd57311;
ROM1[869]<=16'd4779; ROM2[869]<=16'd0; ROM3[869]<=16'd23848; ROM4[869]<=16'd57310;
ROM1[870]<=16'd4774; ROM2[870]<=16'd0; ROM3[870]<=16'd23850; ROM4[870]<=16'd57315;
ROM1[871]<=16'd4778; ROM2[871]<=16'd0; ROM3[871]<=16'd23865; ROM4[871]<=16'd57327;
ROM1[872]<=16'd4780; ROM2[872]<=16'd0; ROM3[872]<=16'd23863; ROM4[872]<=16'd57325;
ROM1[873]<=16'd4780; ROM2[873]<=16'd0; ROM3[873]<=16'd23850; ROM4[873]<=16'd57319;
ROM1[874]<=16'd4807; ROM2[874]<=16'd0; ROM3[874]<=16'd23833; ROM4[874]<=16'd57310;
ROM1[875]<=16'd4843; ROM2[875]<=16'd0; ROM3[875]<=16'd23827; ROM4[875]<=16'd57316;
ROM1[876]<=16'd4846; ROM2[876]<=16'd0; ROM3[876]<=16'd23831; ROM4[876]<=16'd57319;
ROM1[877]<=16'd4809; ROM2[877]<=16'd0; ROM3[877]<=16'd23816; ROM4[877]<=16'd57293;
ROM1[878]<=16'd4798; ROM2[878]<=16'd0; ROM3[878]<=16'd23831; ROM4[878]<=16'd57304;
ROM1[879]<=16'd4794; ROM2[879]<=16'd0; ROM3[879]<=16'd23847; ROM4[879]<=16'd57312;
ROM1[880]<=16'd4791; ROM2[880]<=16'd0; ROM3[880]<=16'd23857; ROM4[880]<=16'd57316;
ROM1[881]<=16'd4816; ROM2[881]<=16'd0; ROM3[881]<=16'd23871; ROM4[881]<=16'd57333;
ROM1[882]<=16'd4851; ROM2[882]<=16'd0; ROM3[882]<=16'd23857; ROM4[882]<=16'd57330;
ROM1[883]<=16'd4882; ROM2[883]<=16'd0; ROM3[883]<=16'd23835; ROM4[883]<=16'd57320;
ROM1[884]<=16'd4891; ROM2[884]<=16'd0; ROM3[884]<=16'd23831; ROM4[884]<=16'd57319;
ROM1[885]<=16'd4892; ROM2[885]<=16'd0; ROM3[885]<=16'd23847; ROM4[885]<=16'd57331;
ROM1[886]<=16'd4900; ROM2[886]<=16'd0; ROM3[886]<=16'd23881; ROM4[886]<=16'd57359;
ROM1[887]<=16'd4898; ROM2[887]<=16'd0; ROM3[887]<=16'd23890; ROM4[887]<=16'd57362;
ROM1[888]<=16'd4883; ROM2[888]<=16'd0; ROM3[888]<=16'd23879; ROM4[888]<=16'd57347;
ROM1[889]<=16'd4911; ROM2[889]<=16'd0; ROM3[889]<=16'd23891; ROM4[889]<=16'd57357;
ROM1[890]<=16'd4944; ROM2[890]<=16'd0; ROM3[890]<=16'd23893; ROM4[890]<=16'd57359;
ROM1[891]<=16'd4969; ROM2[891]<=16'd0; ROM3[891]<=16'd23873; ROM4[891]<=16'd57354;
ROM1[892]<=16'd4997; ROM2[892]<=16'd0; ROM3[892]<=16'd23872; ROM4[892]<=16'd57363;
ROM1[893]<=16'd4993; ROM2[893]<=16'd0; ROM3[893]<=16'd23867; ROM4[893]<=16'd57361;
ROM1[894]<=16'd4974; ROM2[894]<=16'd0; ROM3[894]<=16'd23856; ROM4[894]<=16'd57349;
ROM1[895]<=16'd4968; ROM2[895]<=16'd0; ROM3[895]<=16'd23864; ROM4[895]<=16'd57350;
ROM1[896]<=16'd4959; ROM2[896]<=16'd0; ROM3[896]<=16'd23877; ROM4[896]<=16'd57361;
ROM1[897]<=16'd4954; ROM2[897]<=16'd0; ROM3[897]<=16'd23877; ROM4[897]<=16'd57359;
ROM1[898]<=16'd4961; ROM2[898]<=16'd0; ROM3[898]<=16'd23863; ROM4[898]<=16'd57350;
ROM1[899]<=16'd4987; ROM2[899]<=16'd0; ROM3[899]<=16'd23842; ROM4[899]<=16'd57341;
ROM1[900]<=16'd5025; ROM2[900]<=16'd0; ROM3[900]<=16'd23837; ROM4[900]<=16'd57348;
ROM1[901]<=16'd5021; ROM2[901]<=16'd0; ROM3[901]<=16'd23837; ROM4[901]<=16'd57352;
ROM1[902]<=16'd4994; ROM2[902]<=16'd0; ROM3[902]<=16'd23836; ROM4[902]<=16'd57342;
ROM1[903]<=16'd4977; ROM2[903]<=16'd0; ROM3[903]<=16'd23846; ROM4[903]<=16'd57344;
ROM1[904]<=16'd4966; ROM2[904]<=16'd0; ROM3[904]<=16'd23857; ROM4[904]<=16'd57347;
ROM1[905]<=16'd4951; ROM2[905]<=16'd0; ROM3[905]<=16'd23863; ROM4[905]<=16'd57342;
ROM1[906]<=16'd4948; ROM2[906]<=16'd0; ROM3[906]<=16'd23859; ROM4[906]<=16'd57338;
ROM1[907]<=16'd4980; ROM2[907]<=16'd0; ROM3[907]<=16'd23853; ROM4[907]<=16'd57342;
ROM1[908]<=16'd5006; ROM2[908]<=16'd0; ROM3[908]<=16'd23843; ROM4[908]<=16'd57339;
ROM1[909]<=16'd4998; ROM2[909]<=16'd0; ROM3[909]<=16'd23842; ROM4[909]<=16'd57338;
ROM1[910]<=16'd4993; ROM2[910]<=16'd0; ROM3[910]<=16'd23860; ROM4[910]<=16'd57354;
ROM1[911]<=16'd4986; ROM2[911]<=16'd0; ROM3[911]<=16'd23883; ROM4[911]<=16'd57364;
ROM1[912]<=16'd4964; ROM2[912]<=16'd0; ROM3[912]<=16'd23886; ROM4[912]<=16'd57357;
ROM1[913]<=16'd4936; ROM2[913]<=16'd0; ROM3[913]<=16'd23884; ROM4[913]<=16'd57347;
ROM1[914]<=16'd4931; ROM2[914]<=16'd0; ROM3[914]<=16'd23890; ROM4[914]<=16'd57351;
ROM1[915]<=16'd4946; ROM2[915]<=16'd0; ROM3[915]<=16'd23893; ROM4[915]<=16'd57359;
ROM1[916]<=16'd4976; ROM2[916]<=16'd0; ROM3[916]<=16'd23885; ROM4[916]<=16'd57363;
ROM1[917]<=16'd4993; ROM2[917]<=16'd0; ROM3[917]<=16'd23880; ROM4[917]<=16'd57366;
ROM1[918]<=16'd4995; ROM2[918]<=16'd0; ROM3[918]<=16'd23900; ROM4[918]<=16'd57382;
ROM1[919]<=16'd4948; ROM2[919]<=16'd0; ROM3[919]<=16'd23881; ROM4[919]<=16'd57358;
ROM1[920]<=16'd4890; ROM2[920]<=16'd0; ROM3[920]<=16'd23847; ROM4[920]<=16'd57318;
ROM1[921]<=16'd4869; ROM2[921]<=16'd0; ROM3[921]<=16'd23856; ROM4[921]<=16'd57318;
ROM1[922]<=16'd4850; ROM2[922]<=16'd0; ROM3[922]<=16'd23852; ROM4[922]<=16'd57312;
ROM1[923]<=16'd4873; ROM2[923]<=16'd0; ROM3[923]<=16'd23855; ROM4[923]<=16'd57316;
ROM1[924]<=16'd4927; ROM2[924]<=16'd0; ROM3[924]<=16'd23875; ROM4[924]<=16'd57344;
ROM1[925]<=16'd4934; ROM2[925]<=16'd0; ROM3[925]<=16'd23856; ROM4[925]<=16'd57337;
ROM1[926]<=16'd4899; ROM2[926]<=16'd0; ROM3[926]<=16'd23833; ROM4[926]<=16'd57313;
ROM1[927]<=16'd4880; ROM2[927]<=16'd0; ROM3[927]<=16'd23846; ROM4[927]<=16'd57320;
ROM1[928]<=16'd4870; ROM2[928]<=16'd0; ROM3[928]<=16'd23857; ROM4[928]<=16'd57323;
ROM1[929]<=16'd4830; ROM2[929]<=16'd0; ROM3[929]<=16'd23839; ROM4[929]<=16'd57302;
ROM1[930]<=16'd4814; ROM2[930]<=16'd0; ROM3[930]<=16'd23839; ROM4[930]<=16'd57300;
ROM1[931]<=16'd4812; ROM2[931]<=16'd0; ROM3[931]<=16'd23837; ROM4[931]<=16'd57300;
ROM1[932]<=16'd4826; ROM2[932]<=16'd0; ROM3[932]<=16'd23818; ROM4[932]<=16'd57291;
ROM1[933]<=16'd4867; ROM2[933]<=16'd0; ROM3[933]<=16'd23806; ROM4[933]<=16'd57297;
ROM1[934]<=16'd4865; ROM2[934]<=16'd0; ROM3[934]<=16'd23799; ROM4[934]<=16'd57293;
ROM1[935]<=16'd4839; ROM2[935]<=16'd0; ROM3[935]<=16'd23797; ROM4[935]<=16'd57287;
ROM1[936]<=16'd4824; ROM2[936]<=16'd0; ROM3[936]<=16'd23808; ROM4[936]<=16'd57292;
ROM1[937]<=16'd4814; ROM2[937]<=16'd0; ROM3[937]<=16'd23827; ROM4[937]<=16'd57303;
ROM1[938]<=16'd4794; ROM2[938]<=16'd0; ROM3[938]<=16'd23832; ROM4[938]<=16'd57301;
ROM1[939]<=16'd4790; ROM2[939]<=16'd0; ROM3[939]<=16'd23828; ROM4[939]<=16'd57294;
ROM1[940]<=16'd4810; ROM2[940]<=16'd0; ROM3[940]<=16'd23823; ROM4[940]<=16'd57298;
ROM1[941]<=16'd4846; ROM2[941]<=16'd0; ROM3[941]<=16'd23815; ROM4[941]<=16'd57303;
ROM1[942]<=16'd4859; ROM2[942]<=16'd0; ROM3[942]<=16'd23813; ROM4[942]<=16'd57307;
ROM1[943]<=16'd4856; ROM2[943]<=16'd0; ROM3[943]<=16'd23830; ROM4[943]<=16'd57318;
ROM1[944]<=16'd4867; ROM2[944]<=16'd0; ROM3[944]<=16'd23868; ROM4[944]<=16'd57345;
ROM1[945]<=16'd4846; ROM2[945]<=16'd0; ROM3[945]<=16'd23872; ROM4[945]<=16'd57339;
ROM1[946]<=16'd4806; ROM2[946]<=16'd0; ROM3[946]<=16'd23854; ROM4[946]<=16'd57314;
ROM1[947]<=16'd4784; ROM2[947]<=16'd0; ROM3[947]<=16'd23839; ROM4[947]<=16'd57298;
ROM1[948]<=16'd4778; ROM2[948]<=16'd0; ROM3[948]<=16'd23822; ROM4[948]<=16'd57280;
ROM1[949]<=16'd4817; ROM2[949]<=16'd0; ROM3[949]<=16'd23822; ROM4[949]<=16'd57290;
ROM1[950]<=16'd4857; ROM2[950]<=16'd0; ROM3[950]<=16'd23826; ROM4[950]<=16'd57300;
ROM1[951]<=16'd4850; ROM2[951]<=16'd0; ROM3[951]<=16'd23830; ROM4[951]<=16'd57300;
ROM1[952]<=16'd4829; ROM2[952]<=16'd0; ROM3[952]<=16'd23839; ROM4[952]<=16'd57308;
ROM1[953]<=16'd4840; ROM2[953]<=16'd0; ROM3[953]<=16'd23867; ROM4[953]<=16'd57332;
ROM1[954]<=16'd4825; ROM2[954]<=16'd0; ROM3[954]<=16'd23868; ROM4[954]<=16'd57330;
ROM1[955]<=16'd4787; ROM2[955]<=16'd0; ROM3[955]<=16'd23846; ROM4[955]<=16'd57301;
ROM1[956]<=16'd4784; ROM2[956]<=16'd0; ROM3[956]<=16'd23837; ROM4[956]<=16'd57291;
ROM1[957]<=16'd4785; ROM2[957]<=16'd0; ROM3[957]<=16'd23809; ROM4[957]<=16'd57268;
ROM1[958]<=16'd4816; ROM2[958]<=16'd0; ROM3[958]<=16'd23800; ROM4[958]<=16'd57267;
ROM1[959]<=16'd4835; ROM2[959]<=16'd0; ROM3[959]<=16'd23814; ROM4[959]<=16'd57282;
ROM1[960]<=16'd4816; ROM2[960]<=16'd0; ROM3[960]<=16'd23816; ROM4[960]<=16'd57275;
ROM1[961]<=16'd4809; ROM2[961]<=16'd0; ROM3[961]<=16'd23835; ROM4[961]<=16'd57281;
ROM1[962]<=16'd4812; ROM2[962]<=16'd0; ROM3[962]<=16'd23859; ROM4[962]<=16'd57298;
ROM1[963]<=16'd4806; ROM2[963]<=16'd0; ROM3[963]<=16'd23869; ROM4[963]<=16'd57307;
ROM1[964]<=16'd4795; ROM2[964]<=16'd0; ROM3[964]<=16'd23861; ROM4[964]<=16'd57299;
ROM1[965]<=16'd4801; ROM2[965]<=16'd0; ROM3[965]<=16'd23846; ROM4[965]<=16'd57291;
ROM1[966]<=16'd4845; ROM2[966]<=16'd0; ROM3[966]<=16'd23845; ROM4[966]<=16'd57305;
ROM1[967]<=16'd4859; ROM2[967]<=16'd0; ROM3[967]<=16'd23839; ROM4[967]<=16'd57309;
ROM1[968]<=16'd4838; ROM2[968]<=16'd0; ROM3[968]<=16'd23836; ROM4[968]<=16'd57303;
ROM1[969]<=16'd4822; ROM2[969]<=16'd0; ROM3[969]<=16'd23847; ROM4[969]<=16'd57307;
ROM1[970]<=16'd4815; ROM2[970]<=16'd0; ROM3[970]<=16'd23862; ROM4[970]<=16'd57315;
ROM1[971]<=16'd4812; ROM2[971]<=16'd0; ROM3[971]<=16'd23877; ROM4[971]<=16'd57323;
ROM1[972]<=16'd4799; ROM2[972]<=16'd0; ROM3[972]<=16'd23869; ROM4[972]<=16'd57317;
ROM1[973]<=16'd4806; ROM2[973]<=16'd0; ROM3[973]<=16'd23862; ROM4[973]<=16'd57317;
ROM1[974]<=16'd4821; ROM2[974]<=16'd0; ROM3[974]<=16'd23842; ROM4[974]<=16'd57308;
ROM1[975]<=16'd4827; ROM2[975]<=16'd0; ROM3[975]<=16'd23816; ROM4[975]<=16'd57294;
ROM1[976]<=16'd4833; ROM2[976]<=16'd0; ROM3[976]<=16'd23831; ROM4[976]<=16'd57307;
ROM1[977]<=16'd4813; ROM2[977]<=16'd0; ROM3[977]<=16'd23834; ROM4[977]<=16'd57303;
ROM1[978]<=16'd4788; ROM2[978]<=16'd0; ROM3[978]<=16'd23836; ROM4[978]<=16'd57296;
ROM1[979]<=16'd4780; ROM2[979]<=16'd0; ROM3[979]<=16'd23855; ROM4[979]<=16'd57305;
ROM1[980]<=16'd4777; ROM2[980]<=16'd0; ROM3[980]<=16'd23865; ROM4[980]<=16'd57310;
ROM1[981]<=16'd4780; ROM2[981]<=16'd0; ROM3[981]<=16'd23857; ROM4[981]<=16'd57306;
ROM1[982]<=16'd4797; ROM2[982]<=16'd0; ROM3[982]<=16'd23839; ROM4[982]<=16'd57297;
ROM1[983]<=16'd4829; ROM2[983]<=16'd0; ROM3[983]<=16'd23828; ROM4[983]<=16'd57300;
ROM1[984]<=16'd4841; ROM2[984]<=16'd0; ROM3[984]<=16'd23837; ROM4[984]<=16'd57315;
ROM1[985]<=16'd4820; ROM2[985]<=16'd0; ROM3[985]<=16'd23838; ROM4[985]<=16'd57316;
ROM1[986]<=16'd4781; ROM2[986]<=16'd0; ROM3[986]<=16'd23821; ROM4[986]<=16'd57293;
ROM1[987]<=16'd4774; ROM2[987]<=16'd0; ROM3[987]<=16'd23829; ROM4[987]<=16'd57299;
ROM1[988]<=16'd4770; ROM2[988]<=16'd0; ROM3[988]<=16'd23841; ROM4[988]<=16'd57309;
ROM1[989]<=16'd4766; ROM2[989]<=16'd0; ROM3[989]<=16'd23835; ROM4[989]<=16'd57301;
ROM1[990]<=16'd4799; ROM2[990]<=16'd0; ROM3[990]<=16'd23841; ROM4[990]<=16'd57312;
ROM1[991]<=16'd4830; ROM2[991]<=16'd0; ROM3[991]<=16'd23827; ROM4[991]<=16'd57310;
ROM1[992]<=16'd4821; ROM2[992]<=16'd0; ROM3[992]<=16'd23799; ROM4[992]<=16'd57285;
ROM1[993]<=16'd4819; ROM2[993]<=16'd0; ROM3[993]<=16'd23811; ROM4[993]<=16'd57295;
ROM1[994]<=16'd4811; ROM2[994]<=16'd0; ROM3[994]<=16'd23830; ROM4[994]<=16'd57307;
ROM1[995]<=16'd4781; ROM2[995]<=16'd0; ROM3[995]<=16'd23824; ROM4[995]<=16'd57291;
ROM1[996]<=16'd4769; ROM2[996]<=16'd0; ROM3[996]<=16'd23834; ROM4[996]<=16'd57296;
ROM1[997]<=16'd4762; ROM2[997]<=16'd0; ROM3[997]<=16'd23838; ROM4[997]<=16'd57293;
ROM1[998]<=16'd4758; ROM2[998]<=16'd0; ROM3[998]<=16'd23817; ROM4[998]<=16'd57279;
ROM1[999]<=16'd4786; ROM2[999]<=16'd0; ROM3[999]<=16'd23809; ROM4[999]<=16'd57280;
ROM1[1000]<=16'd4802; ROM2[1000]<=16'd0; ROM3[1000]<=16'd23798; ROM4[1000]<=16'd57275;
ROM1[1001]<=16'd4787; ROM2[1001]<=16'd0; ROM3[1001]<=16'd23794; ROM4[1001]<=16'd57271;
ROM1[1002]<=16'd4772; ROM2[1002]<=16'd0; ROM3[1002]<=16'd23812; ROM4[1002]<=16'd57274;
ROM1[1003]<=16'd4760; ROM2[1003]<=16'd0; ROM3[1003]<=16'd23825; ROM4[1003]<=16'd57276;
ROM1[1004]<=16'd4746; ROM2[1004]<=16'd0; ROM3[1004]<=16'd23824; ROM4[1004]<=16'd57271;
ROM1[1005]<=16'd4732; ROM2[1005]<=16'd0; ROM3[1005]<=16'd23824; ROM4[1005]<=16'd57266;
ROM1[1006]<=16'd4740; ROM2[1006]<=16'd0; ROM3[1006]<=16'd23822; ROM4[1006]<=16'd57267;
ROM1[1007]<=16'd4766; ROM2[1007]<=16'd0; ROM3[1007]<=16'd23806; ROM4[1007]<=16'd57264;
ROM1[1008]<=16'd4797; ROM2[1008]<=16'd0; ROM3[1008]<=16'd23796; ROM4[1008]<=16'd57264;
ROM1[1009]<=16'd4804; ROM2[1009]<=16'd0; ROM3[1009]<=16'd23792; ROM4[1009]<=16'd57267;
ROM1[1010]<=16'd4791; ROM2[1010]<=16'd0; ROM3[1010]<=16'd23796; ROM4[1010]<=16'd57270;
ROM1[1011]<=16'd4779; ROM2[1011]<=16'd0; ROM3[1011]<=16'd23809; ROM4[1011]<=16'd57275;
ROM1[1012]<=16'd4767; ROM2[1012]<=16'd0; ROM3[1012]<=16'd23820; ROM4[1012]<=16'd57283;
ROM1[1013]<=16'd4760; ROM2[1013]<=16'd0; ROM3[1013]<=16'd23832; ROM4[1013]<=16'd57289;
ROM1[1014]<=16'd4775; ROM2[1014]<=16'd0; ROM3[1014]<=16'd23845; ROM4[1014]<=16'd57305;
ROM1[1015]<=16'd4806; ROM2[1015]<=16'd0; ROM3[1015]<=16'd23848; ROM4[1015]<=16'd57316;
ROM1[1016]<=16'd4834; ROM2[1016]<=16'd0; ROM3[1016]<=16'd23837; ROM4[1016]<=16'd57312;
ROM1[1017]<=16'd4842; ROM2[1017]<=16'd0; ROM3[1017]<=16'd23831; ROM4[1017]<=16'd57311;
ROM1[1018]<=16'd4838; ROM2[1018]<=16'd0; ROM3[1018]<=16'd23844; ROM4[1018]<=16'd57319;
ROM1[1019]<=16'd4829; ROM2[1019]<=16'd0; ROM3[1019]<=16'd23862; ROM4[1019]<=16'd57330;
ROM1[1020]<=16'd4801; ROM2[1020]<=16'd0; ROM3[1020]<=16'd23856; ROM4[1020]<=16'd57318;
ROM1[1021]<=16'd4775; ROM2[1021]<=16'd0; ROM3[1021]<=16'd23851; ROM4[1021]<=16'd57308;
ROM1[1022]<=16'd4777; ROM2[1022]<=16'd0; ROM3[1022]<=16'd23855; ROM4[1022]<=16'd57311;
ROM1[1023]<=16'd4791; ROM2[1023]<=16'd0; ROM3[1023]<=16'd23847; ROM4[1023]<=16'd57308;
ROM1[1024]<=16'd4822; ROM2[1024]<=16'd0; ROM3[1024]<=16'd23836; ROM4[1024]<=16'd57303;
ROM1[1025]<=16'd4846; ROM2[1025]<=16'd0; ROM3[1025]<=16'd23827; ROM4[1025]<=16'd57305;
ROM1[1026]<=16'd4815; ROM2[1026]<=16'd0; ROM3[1026]<=16'd23811; ROM4[1026]<=16'd57286;
ROM1[1027]<=16'd4782; ROM2[1027]<=16'd0; ROM3[1027]<=16'd23806; ROM4[1027]<=16'd57271;
ROM1[1028]<=16'd4780; ROM2[1028]<=16'd0; ROM3[1028]<=16'd23821; ROM4[1028]<=16'd57287;
ROM1[1029]<=16'd4776; ROM2[1029]<=16'd0; ROM3[1029]<=16'd23834; ROM4[1029]<=16'd57298;
ROM1[1030]<=16'd4771; ROM2[1030]<=16'd0; ROM3[1030]<=16'd23836; ROM4[1030]<=16'd57299;
ROM1[1031]<=16'd4776; ROM2[1031]<=16'd0; ROM3[1031]<=16'd23828; ROM4[1031]<=16'd57296;
ROM1[1032]<=16'd4793; ROM2[1032]<=16'd0; ROM3[1032]<=16'd23812; ROM4[1032]<=16'd57289;
ROM1[1033]<=16'd4816; ROM2[1033]<=16'd0; ROM3[1033]<=16'd23792; ROM4[1033]<=16'd57284;
ROM1[1034]<=16'd4823; ROM2[1034]<=16'd0; ROM3[1034]<=16'd23792; ROM4[1034]<=16'd57287;
ROM1[1035]<=16'd4804; ROM2[1035]<=16'd0; ROM3[1035]<=16'd23792; ROM4[1035]<=16'd57286;
ROM1[1036]<=16'd4783; ROM2[1036]<=16'd0; ROM3[1036]<=16'd23795; ROM4[1036]<=16'd57280;
ROM1[1037]<=16'd4777; ROM2[1037]<=16'd0; ROM3[1037]<=16'd23807; ROM4[1037]<=16'd57287;
ROM1[1038]<=16'd4771; ROM2[1038]<=16'd0; ROM3[1038]<=16'd23821; ROM4[1038]<=16'd57301;
ROM1[1039]<=16'd4771; ROM2[1039]<=16'd0; ROM3[1039]<=16'd23825; ROM4[1039]<=16'd57302;
ROM1[1040]<=16'd4791; ROM2[1040]<=16'd0; ROM3[1040]<=16'd23821; ROM4[1040]<=16'd57303;
ROM1[1041]<=16'd4813; ROM2[1041]<=16'd0; ROM3[1041]<=16'd23803; ROM4[1041]<=16'd57293;
ROM1[1042]<=16'd4808; ROM2[1042]<=16'd0; ROM3[1042]<=16'd23785; ROM4[1042]<=16'd57274;
ROM1[1043]<=16'd4804; ROM2[1043]<=16'd0; ROM3[1043]<=16'd23799; ROM4[1043]<=16'd57286;
ROM1[1044]<=16'd4787; ROM2[1044]<=16'd0; ROM3[1044]<=16'd23808; ROM4[1044]<=16'd57289;
ROM1[1045]<=16'd4773; ROM2[1045]<=16'd0; ROM3[1045]<=16'd23812; ROM4[1045]<=16'd57289;
ROM1[1046]<=16'd4760; ROM2[1046]<=16'd0; ROM3[1046]<=16'd23820; ROM4[1046]<=16'd57292;
ROM1[1047]<=16'd4749; ROM2[1047]<=16'd0; ROM3[1047]<=16'd23818; ROM4[1047]<=16'd57284;
ROM1[1048]<=16'd4761; ROM2[1048]<=16'd0; ROM3[1048]<=16'd23814; ROM4[1048]<=16'd57284;
ROM1[1049]<=16'd4793; ROM2[1049]<=16'd0; ROM3[1049]<=16'd23804; ROM4[1049]<=16'd57284;
ROM1[1050]<=16'd4812; ROM2[1050]<=16'd0; ROM3[1050]<=16'd23794; ROM4[1050]<=16'd57282;
ROM1[1051]<=16'd4799; ROM2[1051]<=16'd0; ROM3[1051]<=16'd23795; ROM4[1051]<=16'd57280;
ROM1[1052]<=16'd4791; ROM2[1052]<=16'd0; ROM3[1052]<=16'd23819; ROM4[1052]<=16'd57292;
ROM1[1053]<=16'd4785; ROM2[1053]<=16'd0; ROM3[1053]<=16'd23838; ROM4[1053]<=16'd57300;
ROM1[1054]<=16'd4764; ROM2[1054]<=16'd0; ROM3[1054]<=16'd23834; ROM4[1054]<=16'd57292;
ROM1[1055]<=16'd4768; ROM2[1055]<=16'd0; ROM3[1055]<=16'd23846; ROM4[1055]<=16'd57301;
ROM1[1056]<=16'd4788; ROM2[1056]<=16'd0; ROM3[1056]<=16'd23854; ROM4[1056]<=16'd57314;
ROM1[1057]<=16'd4795; ROM2[1057]<=16'd0; ROM3[1057]<=16'd23831; ROM4[1057]<=16'd57299;
ROM1[1058]<=16'd4815; ROM2[1058]<=16'd0; ROM3[1058]<=16'd23809; ROM4[1058]<=16'd57288;
ROM1[1059]<=16'd4820; ROM2[1059]<=16'd0; ROM3[1059]<=16'd23813; ROM4[1059]<=16'd57294;
ROM1[1060]<=16'd4796; ROM2[1060]<=16'd0; ROM3[1060]<=16'd23809; ROM4[1060]<=16'd57285;
ROM1[1061]<=16'd4781; ROM2[1061]<=16'd0; ROM3[1061]<=16'd23822; ROM4[1061]<=16'd57290;
ROM1[1062]<=16'd4769; ROM2[1062]<=16'd0; ROM3[1062]<=16'd23831; ROM4[1062]<=16'd57296;
ROM1[1063]<=16'd4749; ROM2[1063]<=16'd0; ROM3[1063]<=16'd23826; ROM4[1063]<=16'd57286;
ROM1[1064]<=16'd4750; ROM2[1064]<=16'd0; ROM3[1064]<=16'd23823; ROM4[1064]<=16'd57283;
ROM1[1065]<=16'd4763; ROM2[1065]<=16'd0; ROM3[1065]<=16'd23805; ROM4[1065]<=16'd57276;
ROM1[1066]<=16'd4793; ROM2[1066]<=16'd0; ROM3[1066]<=16'd23796; ROM4[1066]<=16'd57274;
ROM1[1067]<=16'd4796; ROM2[1067]<=16'd0; ROM3[1067]<=16'd23787; ROM4[1067]<=16'd57266;
ROM1[1068]<=16'd4777; ROM2[1068]<=16'd0; ROM3[1068]<=16'd23781; ROM4[1068]<=16'd57261;
ROM1[1069]<=16'd4768; ROM2[1069]<=16'd0; ROM3[1069]<=16'd23796; ROM4[1069]<=16'd57270;
ROM1[1070]<=16'd4762; ROM2[1070]<=16'd0; ROM3[1070]<=16'd23815; ROM4[1070]<=16'd57281;
ROM1[1071]<=16'd4750; ROM2[1071]<=16'd0; ROM3[1071]<=16'd23826; ROM4[1071]<=16'd57287;
ROM1[1072]<=16'd4738; ROM2[1072]<=16'd0; ROM3[1072]<=16'd23824; ROM4[1072]<=16'd57280;
ROM1[1073]<=16'd4760; ROM2[1073]<=16'd0; ROM3[1073]<=16'd23830; ROM4[1073]<=16'd57289;
ROM1[1074]<=16'd4814; ROM2[1074]<=16'd0; ROM3[1074]<=16'd23837; ROM4[1074]<=16'd57311;
ROM1[1075]<=16'd4822; ROM2[1075]<=16'd0; ROM3[1075]<=16'd23807; ROM4[1075]<=16'd57295;
ROM1[1076]<=16'd4785; ROM2[1076]<=16'd0; ROM3[1076]<=16'd23782; ROM4[1076]<=16'd57267;
ROM1[1077]<=16'd4761; ROM2[1077]<=16'd0; ROM3[1077]<=16'd23782; ROM4[1077]<=16'd57259;
ROM1[1078]<=16'd4735; ROM2[1078]<=16'd0; ROM3[1078]<=16'd23780; ROM4[1078]<=16'd57250;
ROM1[1079]<=16'd4729; ROM2[1079]<=16'd0; ROM3[1079]<=16'd23796; ROM4[1079]<=16'd57260;
ROM1[1080]<=16'd4744; ROM2[1080]<=16'd0; ROM3[1080]<=16'd23821; ROM4[1080]<=16'd57290;
ROM1[1081]<=16'd4760; ROM2[1081]<=16'd0; ROM3[1081]<=16'd23826; ROM4[1081]<=16'd57301;
ROM1[1082]<=16'd4776; ROM2[1082]<=16'd0; ROM3[1082]<=16'd23805; ROM4[1082]<=16'd57285;
ROM1[1083]<=16'd4802; ROM2[1083]<=16'd0; ROM3[1083]<=16'd23790; ROM4[1083]<=16'd57282;
ROM1[1084]<=16'd4803; ROM2[1084]<=16'd0; ROM3[1084]<=16'd23789; ROM4[1084]<=16'd57282;
ROM1[1085]<=16'd4785; ROM2[1085]<=16'd0; ROM3[1085]<=16'd23794; ROM4[1085]<=16'd57278;
ROM1[1086]<=16'd4783; ROM2[1086]<=16'd0; ROM3[1086]<=16'd23814; ROM4[1086]<=16'd57295;
ROM1[1087]<=16'd4761; ROM2[1087]<=16'd0; ROM3[1087]<=16'd23811; ROM4[1087]<=16'd57285;
ROM1[1088]<=16'd4730; ROM2[1088]<=16'd0; ROM3[1088]<=16'd23801; ROM4[1088]<=16'd57263;
ROM1[1089]<=16'd4728; ROM2[1089]<=16'd0; ROM3[1089]<=16'd23803; ROM4[1089]<=16'd57259;
ROM1[1090]<=16'd4756; ROM2[1090]<=16'd0; ROM3[1090]<=16'd23806; ROM4[1090]<=16'd57268;
ROM1[1091]<=16'd4799; ROM2[1091]<=16'd0; ROM3[1091]<=16'd23802; ROM4[1091]<=16'd57280;
ROM1[1092]<=16'd4804; ROM2[1092]<=16'd0; ROM3[1092]<=16'd23785; ROM4[1092]<=16'd57269;
ROM1[1093]<=16'd4783; ROM2[1093]<=16'd0; ROM3[1093]<=16'd23790; ROM4[1093]<=16'd57267;
ROM1[1094]<=16'd4749; ROM2[1094]<=16'd0; ROM3[1094]<=16'd23792; ROM4[1094]<=16'd57258;
ROM1[1095]<=16'd4731; ROM2[1095]<=16'd0; ROM3[1095]<=16'd23799; ROM4[1095]<=16'd57254;
ROM1[1096]<=16'd4729; ROM2[1096]<=16'd0; ROM3[1096]<=16'd23822; ROM4[1096]<=16'd57270;
ROM1[1097]<=16'd4731; ROM2[1097]<=16'd0; ROM3[1097]<=16'd23825; ROM4[1097]<=16'd57273;
ROM1[1098]<=16'd4740; ROM2[1098]<=16'd0; ROM3[1098]<=16'd23813; ROM4[1098]<=16'd57270;
ROM1[1099]<=16'd4775; ROM2[1099]<=16'd0; ROM3[1099]<=16'd23805; ROM4[1099]<=16'd57275;
ROM1[1100]<=16'd4802; ROM2[1100]<=16'd0; ROM3[1100]<=16'd23797; ROM4[1100]<=16'd57277;
ROM1[1101]<=16'd4788; ROM2[1101]<=16'd0; ROM3[1101]<=16'd23791; ROM4[1101]<=16'd57275;
ROM1[1102]<=16'd4768; ROM2[1102]<=16'd0; ROM3[1102]<=16'd23801; ROM4[1102]<=16'd57275;
ROM1[1103]<=16'd4758; ROM2[1103]<=16'd0; ROM3[1103]<=16'd23818; ROM4[1103]<=16'd57281;
ROM1[1104]<=16'd4759; ROM2[1104]<=16'd0; ROM3[1104]<=16'd23842; ROM4[1104]<=16'd57300;
ROM1[1105]<=16'd4758; ROM2[1105]<=16'd0; ROM3[1105]<=16'd23856; ROM4[1105]<=16'd57307;
ROM1[1106]<=16'd4759; ROM2[1106]<=16'd0; ROM3[1106]<=16'd23842; ROM4[1106]<=16'd57299;
ROM1[1107]<=16'd4784; ROM2[1107]<=16'd0; ROM3[1107]<=16'd23828; ROM4[1107]<=16'd57295;
ROM1[1108]<=16'd4821; ROM2[1108]<=16'd0; ROM3[1108]<=16'd23829; ROM4[1108]<=16'd57300;
ROM1[1109]<=16'd4815; ROM2[1109]<=16'd0; ROM3[1109]<=16'd23818; ROM4[1109]<=16'd57290;
ROM1[1110]<=16'd4791; ROM2[1110]<=16'd0; ROM3[1110]<=16'd23818; ROM4[1110]<=16'd57282;
ROM1[1111]<=16'd4774; ROM2[1111]<=16'd0; ROM3[1111]<=16'd23832; ROM4[1111]<=16'd57287;
ROM1[1112]<=16'd4759; ROM2[1112]<=16'd0; ROM3[1112]<=16'd23835; ROM4[1112]<=16'd57287;
ROM1[1113]<=16'd4741; ROM2[1113]<=16'd0; ROM3[1113]<=16'd23839; ROM4[1113]<=16'd57287;
ROM1[1114]<=16'd4727; ROM2[1114]<=16'd0; ROM3[1114]<=16'd23826; ROM4[1114]<=16'd57274;
ROM1[1115]<=16'd4736; ROM2[1115]<=16'd0; ROM3[1115]<=16'd23811; ROM4[1115]<=16'd57267;
ROM1[1116]<=16'd4766; ROM2[1116]<=16'd0; ROM3[1116]<=16'd23801; ROM4[1116]<=16'd57266;
ROM1[1117]<=16'd4795; ROM2[1117]<=16'd0; ROM3[1117]<=16'd23808; ROM4[1117]<=16'd57281;
ROM1[1118]<=16'd4808; ROM2[1118]<=16'd0; ROM3[1118]<=16'd23835; ROM4[1118]<=16'd57306;
ROM1[1119]<=16'd4778; ROM2[1119]<=16'd0; ROM3[1119]<=16'd23830; ROM4[1119]<=16'd57294;
ROM1[1120]<=16'd4746; ROM2[1120]<=16'd0; ROM3[1120]<=16'd23818; ROM4[1120]<=16'd57282;
ROM1[1121]<=16'd4733; ROM2[1121]<=16'd0; ROM3[1121]<=16'd23826; ROM4[1121]<=16'd57281;
ROM1[1122]<=16'd4734; ROM2[1122]<=16'd0; ROM3[1122]<=16'd23829; ROM4[1122]<=16'd57282;
ROM1[1123]<=16'd4759; ROM2[1123]<=16'd0; ROM3[1123]<=16'd23830; ROM4[1123]<=16'd57289;
ROM1[1124]<=16'd4792; ROM2[1124]<=16'd0; ROM3[1124]<=16'd23827; ROM4[1124]<=16'd57294;
ROM1[1125]<=16'd4814; ROM2[1125]<=16'd0; ROM3[1125]<=16'd23818; ROM4[1125]<=16'd57301;
ROM1[1126]<=16'd4802; ROM2[1126]<=16'd0; ROM3[1126]<=16'd23809; ROM4[1126]<=16'd57290;
ROM1[1127]<=16'd4771; ROM2[1127]<=16'd0; ROM3[1127]<=16'd23800; ROM4[1127]<=16'd57278;
ROM1[1128]<=16'd4754; ROM2[1128]<=16'd0; ROM3[1128]<=16'd23798; ROM4[1128]<=16'd57273;
ROM1[1129]<=16'd4735; ROM2[1129]<=16'd0; ROM3[1129]<=16'd23799; ROM4[1129]<=16'd57265;
ROM1[1130]<=16'd4727; ROM2[1130]<=16'd0; ROM3[1130]<=16'd23805; ROM4[1130]<=16'd57269;
ROM1[1131]<=16'd4744; ROM2[1131]<=16'd0; ROM3[1131]<=16'd23813; ROM4[1131]<=16'd57277;
ROM1[1132]<=16'd4774; ROM2[1132]<=16'd0; ROM3[1132]<=16'd23811; ROM4[1132]<=16'd57283;
ROM1[1133]<=16'd4800; ROM2[1133]<=16'd0; ROM3[1133]<=16'd23798; ROM4[1133]<=16'd57282;
ROM1[1134]<=16'd4800; ROM2[1134]<=16'd0; ROM3[1134]<=16'd23796; ROM4[1134]<=16'd57282;
ROM1[1135]<=16'd4803; ROM2[1135]<=16'd0; ROM3[1135]<=16'd23821; ROM4[1135]<=16'd57302;
ROM1[1136]<=16'd4790; ROM2[1136]<=16'd0; ROM3[1136]<=16'd23838; ROM4[1136]<=16'd57310;
ROM1[1137]<=16'd4762; ROM2[1137]<=16'd0; ROM3[1137]<=16'd23828; ROM4[1137]<=16'd57294;
ROM1[1138]<=16'd4743; ROM2[1138]<=16'd0; ROM3[1138]<=16'd23822; ROM4[1138]<=16'd57288;
ROM1[1139]<=16'd4732; ROM2[1139]<=16'd0; ROM3[1139]<=16'd23815; ROM4[1139]<=16'd57281;
ROM1[1140]<=16'd4743; ROM2[1140]<=16'd0; ROM3[1140]<=16'd23798; ROM4[1140]<=16'd57270;
ROM1[1141]<=16'd4778; ROM2[1141]<=16'd0; ROM3[1141]<=16'd23789; ROM4[1141]<=16'd57274;
ROM1[1142]<=16'd4791; ROM2[1142]<=16'd0; ROM3[1142]<=16'd23794; ROM4[1142]<=16'd57278;
ROM1[1143]<=16'd4779; ROM2[1143]<=16'd0; ROM3[1143]<=16'd23800; ROM4[1143]<=16'd57276;
ROM1[1144]<=16'd4766; ROM2[1144]<=16'd0; ROM3[1144]<=16'd23816; ROM4[1144]<=16'd57287;
ROM1[1145]<=16'd4758; ROM2[1145]<=16'd0; ROM3[1145]<=16'd23837; ROM4[1145]<=16'd57300;
ROM1[1146]<=16'd4738; ROM2[1146]<=16'd0; ROM3[1146]<=16'd23844; ROM4[1146]<=16'd57302;
ROM1[1147]<=16'd4732; ROM2[1147]<=16'd0; ROM3[1147]<=16'd23848; ROM4[1147]<=16'd57301;
ROM1[1148]<=16'd4743; ROM2[1148]<=16'd0; ROM3[1148]<=16'd23840; ROM4[1148]<=16'd57297;
ROM1[1149]<=16'd4773; ROM2[1149]<=16'd0; ROM3[1149]<=16'd23826; ROM4[1149]<=16'd57296;
ROM1[1150]<=16'd4804; ROM2[1150]<=16'd0; ROM3[1150]<=16'd23825; ROM4[1150]<=16'd57305;
ROM1[1151]<=16'd4799; ROM2[1151]<=16'd0; ROM3[1151]<=16'd23827; ROM4[1151]<=16'd57307;
ROM1[1152]<=16'd4778; ROM2[1152]<=16'd0; ROM3[1152]<=16'd23827; ROM4[1152]<=16'd57301;
ROM1[1153]<=16'd4763; ROM2[1153]<=16'd0; ROM3[1153]<=16'd23830; ROM4[1153]<=16'd57296;
ROM1[1154]<=16'd4749; ROM2[1154]<=16'd0; ROM3[1154]<=16'd23832; ROM4[1154]<=16'd57290;
ROM1[1155]<=16'd4738; ROM2[1155]<=16'd0; ROM3[1155]<=16'd23833; ROM4[1155]<=16'd57289;
ROM1[1156]<=16'd4751; ROM2[1156]<=16'd0; ROM3[1156]<=16'd23835; ROM4[1156]<=16'd57297;
ROM1[1157]<=16'd4780; ROM2[1157]<=16'd0; ROM3[1157]<=16'd23833; ROM4[1157]<=16'd57302;
ROM1[1158]<=16'd4807; ROM2[1158]<=16'd0; ROM3[1158]<=16'd23825; ROM4[1158]<=16'd57301;
ROM1[1159]<=16'd4813; ROM2[1159]<=16'd0; ROM3[1159]<=16'd23827; ROM4[1159]<=16'd57304;
ROM1[1160]<=16'd4811; ROM2[1160]<=16'd0; ROM3[1160]<=16'd23844; ROM4[1160]<=16'd57319;
ROM1[1161]<=16'd4786; ROM2[1161]<=16'd0; ROM3[1161]<=16'd23846; ROM4[1161]<=16'd57315;
ROM1[1162]<=16'd4759; ROM2[1162]<=16'd0; ROM3[1162]<=16'd23838; ROM4[1162]<=16'd57302;
ROM1[1163]<=16'd4747; ROM2[1163]<=16'd0; ROM3[1163]<=16'd23850; ROM4[1163]<=16'd57307;
ROM1[1164]<=16'd4747; ROM2[1164]<=16'd0; ROM3[1164]<=16'd23849; ROM4[1164]<=16'd57304;
ROM1[1165]<=16'd4770; ROM2[1165]<=16'd0; ROM3[1165]<=16'd23845; ROM4[1165]<=16'd57309;
ROM1[1166]<=16'd4814; ROM2[1166]<=16'd0; ROM3[1166]<=16'd23848; ROM4[1166]<=16'd57321;
ROM1[1167]<=16'd4825; ROM2[1167]<=16'd0; ROM3[1167]<=16'd23841; ROM4[1167]<=16'd57321;
ROM1[1168]<=16'd4797; ROM2[1168]<=16'd0; ROM3[1168]<=16'd23830; ROM4[1168]<=16'd57307;
ROM1[1169]<=16'd4774; ROM2[1169]<=16'd0; ROM3[1169]<=16'd23833; ROM4[1169]<=16'd57299;
ROM1[1170]<=16'd4759; ROM2[1170]<=16'd0; ROM3[1170]<=16'd23834; ROM4[1170]<=16'd57297;
ROM1[1171]<=16'd4745; ROM2[1171]<=16'd0; ROM3[1171]<=16'd23840; ROM4[1171]<=16'd57296;
ROM1[1172]<=16'd4747; ROM2[1172]<=16'd0; ROM3[1172]<=16'd23849; ROM4[1172]<=16'd57304;
ROM1[1173]<=16'd4759; ROM2[1173]<=16'd0; ROM3[1173]<=16'd23843; ROM4[1173]<=16'd57302;
ROM1[1174]<=16'd4790; ROM2[1174]<=16'd0; ROM3[1174]<=16'd23829; ROM4[1174]<=16'd57301;
ROM1[1175]<=16'd4813; ROM2[1175]<=16'd0; ROM3[1175]<=16'd23823; ROM4[1175]<=16'd57305;
ROM1[1176]<=16'd4800; ROM2[1176]<=16'd0; ROM3[1176]<=16'd23825; ROM4[1176]<=16'd57302;
ROM1[1177]<=16'd4785; ROM2[1177]<=16'd0; ROM3[1177]<=16'd23830; ROM4[1177]<=16'd57306;
ROM1[1178]<=16'd4778; ROM2[1178]<=16'd0; ROM3[1178]<=16'd23843; ROM4[1178]<=16'd57316;
ROM1[1179]<=16'd4783; ROM2[1179]<=16'd0; ROM3[1179]<=16'd23865; ROM4[1179]<=16'd57332;
ROM1[1180]<=16'd4769; ROM2[1180]<=16'd0; ROM3[1180]<=16'd23860; ROM4[1180]<=16'd57324;
ROM1[1181]<=16'd4745; ROM2[1181]<=16'd0; ROM3[1181]<=16'd23828; ROM4[1181]<=16'd57293;
ROM1[1182]<=16'd4760; ROM2[1182]<=16'd0; ROM3[1182]<=16'd23806; ROM4[1182]<=16'd57278;
ROM1[1183]<=16'd4776; ROM2[1183]<=16'd0; ROM3[1183]<=16'd23784; ROM4[1183]<=16'd57267;
ROM1[1184]<=16'd4775; ROM2[1184]<=16'd0; ROM3[1184]<=16'd23787; ROM4[1184]<=16'd57270;
ROM1[1185]<=16'd4779; ROM2[1185]<=16'd0; ROM3[1185]<=16'd23811; ROM4[1185]<=16'd57292;
ROM1[1186]<=16'd4757; ROM2[1186]<=16'd0; ROM3[1186]<=16'd23819; ROM4[1186]<=16'd57287;
ROM1[1187]<=16'd4729; ROM2[1187]<=16'd0; ROM3[1187]<=16'd23804; ROM4[1187]<=16'd57268;
ROM1[1188]<=16'd4719; ROM2[1188]<=16'd0; ROM3[1188]<=16'd23804; ROM4[1188]<=16'd57267;
ROM1[1189]<=16'd4734; ROM2[1189]<=16'd0; ROM3[1189]<=16'd23815; ROM4[1189]<=16'd57275;
ROM1[1190]<=16'd4757; ROM2[1190]<=16'd0; ROM3[1190]<=16'd23806; ROM4[1190]<=16'd57276;
ROM1[1191]<=16'd4788; ROM2[1191]<=16'd0; ROM3[1191]<=16'd23798; ROM4[1191]<=16'd57276;
ROM1[1192]<=16'd4813; ROM2[1192]<=16'd0; ROM3[1192]<=16'd23814; ROM4[1192]<=16'd57291;
ROM1[1193]<=16'd4825; ROM2[1193]<=16'd0; ROM3[1193]<=16'd23847; ROM4[1193]<=16'd57318;
ROM1[1194]<=16'd4793; ROM2[1194]<=16'd0; ROM3[1194]<=16'd23840; ROM4[1194]<=16'd57308;
ROM1[1195]<=16'd4756; ROM2[1195]<=16'd0; ROM3[1195]<=16'd23821; ROM4[1195]<=16'd57282;
ROM1[1196]<=16'd4735; ROM2[1196]<=16'd0; ROM3[1196]<=16'd23818; ROM4[1196]<=16'd57275;
ROM1[1197]<=16'd4726; ROM2[1197]<=16'd0; ROM3[1197]<=16'd23813; ROM4[1197]<=16'd57267;
ROM1[1198]<=16'd4761; ROM2[1198]<=16'd0; ROM3[1198]<=16'd23827; ROM4[1198]<=16'd57284;
ROM1[1199]<=16'd4819; ROM2[1199]<=16'd0; ROM3[1199]<=16'd23845; ROM4[1199]<=16'd57313;
ROM1[1200]<=16'd4852; ROM2[1200]<=16'd0; ROM3[1200]<=16'd23849; ROM4[1200]<=16'd57326;
ROM1[1201]<=16'd4825; ROM2[1201]<=16'd0; ROM3[1201]<=16'd23837; ROM4[1201]<=16'd57311;
ROM1[1202]<=16'd4793; ROM2[1202]<=16'd0; ROM3[1202]<=16'd23830; ROM4[1202]<=16'd57299;
ROM1[1203]<=16'd4775; ROM2[1203]<=16'd0; ROM3[1203]<=16'd23834; ROM4[1203]<=16'd57301;
ROM1[1204]<=16'd4756; ROM2[1204]<=16'd0; ROM3[1204]<=16'd23836; ROM4[1204]<=16'd57298;
ROM1[1205]<=16'd4760; ROM2[1205]<=16'd0; ROM3[1205]<=16'd23848; ROM4[1205]<=16'd57304;
ROM1[1206]<=16'd4775; ROM2[1206]<=16'd0; ROM3[1206]<=16'd23847; ROM4[1206]<=16'd57305;
ROM1[1207]<=16'd4786; ROM2[1207]<=16'd0; ROM3[1207]<=16'd23818; ROM4[1207]<=16'd57288;
ROM1[1208]<=16'd4806; ROM2[1208]<=16'd0; ROM3[1208]<=16'd23802; ROM4[1208]<=16'd57281;
ROM1[1209]<=16'd4802; ROM2[1209]<=16'd0; ROM3[1209]<=16'd23801; ROM4[1209]<=16'd57279;
ROM1[1210]<=16'd4789; ROM2[1210]<=16'd0; ROM3[1210]<=16'd23819; ROM4[1210]<=16'd57289;
ROM1[1211]<=16'd4777; ROM2[1211]<=16'd0; ROM3[1211]<=16'd23835; ROM4[1211]<=16'd57296;
ROM1[1212]<=16'd4751; ROM2[1212]<=16'd0; ROM3[1212]<=16'd23822; ROM4[1212]<=16'd57281;
ROM1[1213]<=16'd4726; ROM2[1213]<=16'd0; ROM3[1213]<=16'd23815; ROM4[1213]<=16'd57271;
ROM1[1214]<=16'd4736; ROM2[1214]<=16'd0; ROM3[1214]<=16'd23822; ROM4[1214]<=16'd57278;
ROM1[1215]<=16'd4776; ROM2[1215]<=16'd0; ROM3[1215]<=16'd23831; ROM4[1215]<=16'd57293;
ROM1[1216]<=16'd4808; ROM2[1216]<=16'd0; ROM3[1216]<=16'd23824; ROM4[1216]<=16'd57296;
ROM1[1217]<=16'd4803; ROM2[1217]<=16'd0; ROM3[1217]<=16'd23807; ROM4[1217]<=16'd57285;
ROM1[1218]<=16'd4795; ROM2[1218]<=16'd0; ROM3[1218]<=16'd23820; ROM4[1218]<=16'd57294;
ROM1[1219]<=16'd4787; ROM2[1219]<=16'd0; ROM3[1219]<=16'd23838; ROM4[1219]<=16'd57307;
ROM1[1220]<=16'd4766; ROM2[1220]<=16'd0; ROM3[1220]<=16'd23829; ROM4[1220]<=16'd57296;
ROM1[1221]<=16'd4742; ROM2[1221]<=16'd0; ROM3[1221]<=16'd23824; ROM4[1221]<=16'd57288;
ROM1[1222]<=16'd4732; ROM2[1222]<=16'd0; ROM3[1222]<=16'd23819; ROM4[1222]<=16'd57282;
ROM1[1223]<=16'd4746; ROM2[1223]<=16'd0; ROM3[1223]<=16'd23818; ROM4[1223]<=16'd57285;
ROM1[1224]<=16'd4793; ROM2[1224]<=16'd0; ROM3[1224]<=16'd23823; ROM4[1224]<=16'd57301;
ROM1[1225]<=16'd4829; ROM2[1225]<=16'd0; ROM3[1225]<=16'd23821; ROM4[1225]<=16'd57309;
ROM1[1226]<=16'd4810; ROM2[1226]<=16'd0; ROM3[1226]<=16'd23811; ROM4[1226]<=16'd57298;
ROM1[1227]<=16'd4781; ROM2[1227]<=16'd0; ROM3[1227]<=16'd23804; ROM4[1227]<=16'd57287;
ROM1[1228]<=16'd4769; ROM2[1228]<=16'd0; ROM3[1228]<=16'd23812; ROM4[1228]<=16'd57288;
ROM1[1229]<=16'd4776; ROM2[1229]<=16'd0; ROM3[1229]<=16'd23837; ROM4[1229]<=16'd57304;
ROM1[1230]<=16'd4778; ROM2[1230]<=16'd0; ROM3[1230]<=16'd23851; ROM4[1230]<=16'd57314;
ROM1[1231]<=16'd4767; ROM2[1231]<=16'd0; ROM3[1231]<=16'd23835; ROM4[1231]<=16'd57295;
ROM1[1232]<=16'd4791; ROM2[1232]<=16'd0; ROM3[1232]<=16'd23822; ROM4[1232]<=16'd57293;
ROM1[1233]<=16'd4818; ROM2[1233]<=16'd0; ROM3[1233]<=16'd23810; ROM4[1233]<=16'd57294;
ROM1[1234]<=16'd4807; ROM2[1234]<=16'd0; ROM3[1234]<=16'd23802; ROM4[1234]<=16'd57287;
ROM1[1235]<=16'd4799; ROM2[1235]<=16'd0; ROM3[1235]<=16'd23815; ROM4[1235]<=16'd57293;
ROM1[1236]<=16'd4792; ROM2[1236]<=16'd0; ROM3[1236]<=16'd23835; ROM4[1236]<=16'd57303;
ROM1[1237]<=16'd4775; ROM2[1237]<=16'd0; ROM3[1237]<=16'd23839; ROM4[1237]<=16'd57300;
ROM1[1238]<=16'd4759; ROM2[1238]<=16'd0; ROM3[1238]<=16'd23844; ROM4[1238]<=16'd57300;
ROM1[1239]<=16'd4762; ROM2[1239]<=16'd0; ROM3[1239]<=16'd23844; ROM4[1239]<=16'd57299;
ROM1[1240]<=16'd4777; ROM2[1240]<=16'd0; ROM3[1240]<=16'd23834; ROM4[1240]<=16'd57293;
ROM1[1241]<=16'd4811; ROM2[1241]<=16'd0; ROM3[1241]<=16'd23823; ROM4[1241]<=16'd57296;
ROM1[1242]<=16'd4825; ROM2[1242]<=16'd0; ROM3[1242]<=16'd23817; ROM4[1242]<=16'd57296;
ROM1[1243]<=16'd4815; ROM2[1243]<=16'd0; ROM3[1243]<=16'd23825; ROM4[1243]<=16'd57298;
ROM1[1244]<=16'd4805; ROM2[1244]<=16'd0; ROM3[1244]<=16'd23840; ROM4[1244]<=16'd57306;
ROM1[1245]<=16'd4797; ROM2[1245]<=16'd0; ROM3[1245]<=16'd23849; ROM4[1245]<=16'd57308;
ROM1[1246]<=16'd4788; ROM2[1246]<=16'd0; ROM3[1246]<=16'd23860; ROM4[1246]<=16'd57315;
ROM1[1247]<=16'd4792; ROM2[1247]<=16'd0; ROM3[1247]<=16'd23867; ROM4[1247]<=16'd57321;
ROM1[1248]<=16'd4801; ROM2[1248]<=16'd0; ROM3[1248]<=16'd23859; ROM4[1248]<=16'd57315;
ROM1[1249]<=16'd4808; ROM2[1249]<=16'd0; ROM3[1249]<=16'd23832; ROM4[1249]<=16'd57294;
ROM1[1250]<=16'd4848; ROM2[1250]<=16'd0; ROM3[1250]<=16'd23836; ROM4[1250]<=16'd57309;
ROM1[1251]<=16'd4869; ROM2[1251]<=16'd0; ROM3[1251]<=16'd23862; ROM4[1251]<=16'd57334;
ROM1[1252]<=16'd4822; ROM2[1252]<=16'd0; ROM3[1252]<=16'd23837; ROM4[1252]<=16'd57306;
ROM1[1253]<=16'd4782; ROM2[1253]<=16'd0; ROM3[1253]<=16'd23824; ROM4[1253]<=16'd57286;
ROM1[1254]<=16'd4756; ROM2[1254]<=16'd0; ROM3[1254]<=16'd23819; ROM4[1254]<=16'd57280;
ROM1[1255]<=16'd4730; ROM2[1255]<=16'd0; ROM3[1255]<=16'd23804; ROM4[1255]<=16'd57263;
ROM1[1256]<=16'd4755; ROM2[1256]<=16'd0; ROM3[1256]<=16'd23820; ROM4[1256]<=16'd57281;
ROM1[1257]<=16'd4798; ROM2[1257]<=16'd0; ROM3[1257]<=16'd23826; ROM4[1257]<=16'd57299;
ROM1[1258]<=16'd4822; ROM2[1258]<=16'd0; ROM3[1258]<=16'd23816; ROM4[1258]<=16'd57295;
ROM1[1259]<=16'd4816; ROM2[1259]<=16'd0; ROM3[1259]<=16'd23813; ROM4[1259]<=16'd57292;
ROM1[1260]<=16'd4802; ROM2[1260]<=16'd0; ROM3[1260]<=16'd23819; ROM4[1260]<=16'd57293;
ROM1[1261]<=16'd4787; ROM2[1261]<=16'd0; ROM3[1261]<=16'd23823; ROM4[1261]<=16'd57291;
ROM1[1262]<=16'd4761; ROM2[1262]<=16'd0; ROM3[1262]<=16'd23817; ROM4[1262]<=16'd57280;
ROM1[1263]<=16'd4736; ROM2[1263]<=16'd0; ROM3[1263]<=16'd23819; ROM4[1263]<=16'd57271;
ROM1[1264]<=16'd4730; ROM2[1264]<=16'd0; ROM3[1264]<=16'd23817; ROM4[1264]<=16'd57270;
ROM1[1265]<=16'd4751; ROM2[1265]<=16'd0; ROM3[1265]<=16'd23812; ROM4[1265]<=16'd57269;
ROM1[1266]<=16'd4788; ROM2[1266]<=16'd0; ROM3[1266]<=16'd23805; ROM4[1266]<=16'd57268;
ROM1[1267]<=16'd4782; ROM2[1267]<=16'd0; ROM3[1267]<=16'd23782; ROM4[1267]<=16'd57253;
ROM1[1268]<=16'd4751; ROM2[1268]<=16'd0; ROM3[1268]<=16'd23766; ROM4[1268]<=16'd57237;
ROM1[1269]<=16'd4730; ROM2[1269]<=16'd0; ROM3[1269]<=16'd23769; ROM4[1269]<=16'd57235;
ROM1[1270]<=16'd4719; ROM2[1270]<=16'd0; ROM3[1270]<=16'd23778; ROM4[1270]<=16'd57242;
ROM1[1271]<=16'd4712; ROM2[1271]<=16'd0; ROM3[1271]<=16'd23792; ROM4[1271]<=16'd57249;
ROM1[1272]<=16'd4712; ROM2[1272]<=16'd0; ROM3[1272]<=16'd23796; ROM4[1272]<=16'd57253;
ROM1[1273]<=16'd4737; ROM2[1273]<=16'd0; ROM3[1273]<=16'd23800; ROM4[1273]<=16'd57261;
ROM1[1274]<=16'd4777; ROM2[1274]<=16'd0; ROM3[1274]<=16'd23796; ROM4[1274]<=16'd57264;
ROM1[1275]<=16'd4792; ROM2[1275]<=16'd0; ROM3[1275]<=16'd23781; ROM4[1275]<=16'd57262;
ROM1[1276]<=16'd4795; ROM2[1276]<=16'd0; ROM3[1276]<=16'd23799; ROM4[1276]<=16'd57275;
ROM1[1277]<=16'd4784; ROM2[1277]<=16'd0; ROM3[1277]<=16'd23820; ROM4[1277]<=16'd57288;
ROM1[1278]<=16'd4762; ROM2[1278]<=16'd0; ROM3[1278]<=16'd23825; ROM4[1278]<=16'd57285;
ROM1[1279]<=16'd4753; ROM2[1279]<=16'd0; ROM3[1279]<=16'd23835; ROM4[1279]<=16'd57289;
ROM1[1280]<=16'd4747; ROM2[1280]<=16'd0; ROM3[1280]<=16'd23839; ROM4[1280]<=16'd57290;
ROM1[1281]<=16'd4758; ROM2[1281]<=16'd0; ROM3[1281]<=16'd23838; ROM4[1281]<=16'd57290;
ROM1[1282]<=16'd4785; ROM2[1282]<=16'd0; ROM3[1282]<=16'd23828; ROM4[1282]<=16'd57292;
ROM1[1283]<=16'd4819; ROM2[1283]<=16'd0; ROM3[1283]<=16'd23822; ROM4[1283]<=16'd57299;
ROM1[1284]<=16'd4823; ROM2[1284]<=16'd0; ROM3[1284]<=16'd23830; ROM4[1284]<=16'd57307;
ROM1[1285]<=16'd4812; ROM2[1285]<=16'd0; ROM3[1285]<=16'd23843; ROM4[1285]<=16'd57313;
ROM1[1286]<=16'd4803; ROM2[1286]<=16'd0; ROM3[1286]<=16'd23855; ROM4[1286]<=16'd57314;
ROM1[1287]<=16'd4785; ROM2[1287]<=16'd0; ROM3[1287]<=16'd23856; ROM4[1287]<=16'd57311;
ROM1[1288]<=16'd4773; ROM2[1288]<=16'd0; ROM3[1288]<=16'd23863; ROM4[1288]<=16'd57315;
ROM1[1289]<=16'd4775; ROM2[1289]<=16'd0; ROM3[1289]<=16'd23859; ROM4[1289]<=16'd57315;
ROM1[1290]<=16'd4783; ROM2[1290]<=16'd0; ROM3[1290]<=16'd23840; ROM4[1290]<=16'd57305;
ROM1[1291]<=16'd4820; ROM2[1291]<=16'd0; ROM3[1291]<=16'd23836; ROM4[1291]<=16'd57308;
ROM1[1292]<=16'd4845; ROM2[1292]<=16'd0; ROM3[1292]<=16'd23840; ROM4[1292]<=16'd57316;
ROM1[1293]<=16'd4839; ROM2[1293]<=16'd0; ROM3[1293]<=16'd23850; ROM4[1293]<=16'd57321;
ROM1[1294]<=16'd4816; ROM2[1294]<=16'd0; ROM3[1294]<=16'd23857; ROM4[1294]<=16'd57317;
ROM1[1295]<=16'd4794; ROM2[1295]<=16'd0; ROM3[1295]<=16'd23855; ROM4[1295]<=16'd57307;
ROM1[1296]<=16'd4786; ROM2[1296]<=16'd0; ROM3[1296]<=16'd23867; ROM4[1296]<=16'd57312;
ROM1[1297]<=16'd4778; ROM2[1297]<=16'd0; ROM3[1297]<=16'd23868; ROM4[1297]<=16'd57309;
ROM1[1298]<=16'd4790; ROM2[1298]<=16'd0; ROM3[1298]<=16'd23857; ROM4[1298]<=16'd57304;
ROM1[1299]<=16'd4818; ROM2[1299]<=16'd0; ROM3[1299]<=16'd23833; ROM4[1299]<=16'd57295;
ROM1[1300]<=16'd4816; ROM2[1300]<=16'd0; ROM3[1300]<=16'd23802; ROM4[1300]<=16'd57277;
ROM1[1301]<=16'd4803; ROM2[1301]<=16'd0; ROM3[1301]<=16'd23797; ROM4[1301]<=16'd57274;
ROM1[1302]<=16'd4790; ROM2[1302]<=16'd0; ROM3[1302]<=16'd23809; ROM4[1302]<=16'd57279;
ROM1[1303]<=16'd4782; ROM2[1303]<=16'd0; ROM3[1303]<=16'd23825; ROM4[1303]<=16'd57286;
ROM1[1304]<=16'd4782; ROM2[1304]<=16'd0; ROM3[1304]<=16'd23839; ROM4[1304]<=16'd57296;
ROM1[1305]<=16'd4779; ROM2[1305]<=16'd0; ROM3[1305]<=16'd23845; ROM4[1305]<=16'd57298;
ROM1[1306]<=16'd4781; ROM2[1306]<=16'd0; ROM3[1306]<=16'd23833; ROM4[1306]<=16'd57290;
ROM1[1307]<=16'd4799; ROM2[1307]<=16'd0; ROM3[1307]<=16'd23818; ROM4[1307]<=16'd57286;
ROM1[1308]<=16'd4824; ROM2[1308]<=16'd0; ROM3[1308]<=16'd23803; ROM4[1308]<=16'd57281;
ROM1[1309]<=16'd4813; ROM2[1309]<=16'd0; ROM3[1309]<=16'd23794; ROM4[1309]<=16'd57277;
ROM1[1310]<=16'd4807; ROM2[1310]<=16'd0; ROM3[1310]<=16'd23812; ROM4[1310]<=16'd57290;
ROM1[1311]<=16'd4808; ROM2[1311]<=16'd0; ROM3[1311]<=16'd23834; ROM4[1311]<=16'd57302;
ROM1[1312]<=16'd4803; ROM2[1312]<=16'd0; ROM3[1312]<=16'd23852; ROM4[1312]<=16'd57315;
ROM1[1313]<=16'd4800; ROM2[1313]<=16'd0; ROM3[1313]<=16'd23864; ROM4[1313]<=16'd57324;
ROM1[1314]<=16'd4806; ROM2[1314]<=16'd0; ROM3[1314]<=16'd23871; ROM4[1314]<=16'd57328;
ROM1[1315]<=16'd4811; ROM2[1315]<=16'd0; ROM3[1315]<=16'd23847; ROM4[1315]<=16'd57312;
ROM1[1316]<=16'd4810; ROM2[1316]<=16'd0; ROM3[1316]<=16'd23801; ROM4[1316]<=16'd57280;
ROM1[1317]<=16'd4814; ROM2[1317]<=16'd0; ROM3[1317]<=16'd23793; ROM4[1317]<=16'd57277;
ROM1[1318]<=16'd4807; ROM2[1318]<=16'd0; ROM3[1318]<=16'd23797; ROM4[1318]<=16'd57277;
ROM1[1319]<=16'd4799; ROM2[1319]<=16'd0; ROM3[1319]<=16'd23808; ROM4[1319]<=16'd57284;
ROM1[1320]<=16'd4802; ROM2[1320]<=16'd0; ROM3[1320]<=16'd23834; ROM4[1320]<=16'd57301;
ROM1[1321]<=16'd4778; ROM2[1321]<=16'd0; ROM3[1321]<=16'd23836; ROM4[1321]<=16'd57293;
ROM1[1322]<=16'd4762; ROM2[1322]<=16'd0; ROM3[1322]<=16'd23826; ROM4[1322]<=16'd57290;
ROM1[1323]<=16'd4776; ROM2[1323]<=16'd0; ROM3[1323]<=16'd23825; ROM4[1323]<=16'd57293;
ROM1[1324]<=16'd4816; ROM2[1324]<=16'd0; ROM3[1324]<=16'd23820; ROM4[1324]<=16'd57299;
ROM1[1325]<=16'd4851; ROM2[1325]<=16'd0; ROM3[1325]<=16'd23821; ROM4[1325]<=16'd57312;
ROM1[1326]<=16'd4853; ROM2[1326]<=16'd0; ROM3[1326]<=16'd23831; ROM4[1326]<=16'd57319;
ROM1[1327]<=16'd4831; ROM2[1327]<=16'd0; ROM3[1327]<=16'd23838; ROM4[1327]<=16'd57318;
ROM1[1328]<=16'd4808; ROM2[1328]<=16'd0; ROM3[1328]<=16'd23837; ROM4[1328]<=16'd57310;
ROM1[1329]<=16'd4788; ROM2[1329]<=16'd0; ROM3[1329]<=16'd23840; ROM4[1329]<=16'd57304;
ROM1[1330]<=16'd4781; ROM2[1330]<=16'd0; ROM3[1330]<=16'd23846; ROM4[1330]<=16'd57304;
ROM1[1331]<=16'd4793; ROM2[1331]<=16'd0; ROM3[1331]<=16'd23845; ROM4[1331]<=16'd57301;
ROM1[1332]<=16'd4819; ROM2[1332]<=16'd0; ROM3[1332]<=16'd23839; ROM4[1332]<=16'd57302;
ROM1[1333]<=16'd4841; ROM2[1333]<=16'd0; ROM3[1333]<=16'd23829; ROM4[1333]<=16'd57300;
ROM1[1334]<=16'd4834; ROM2[1334]<=16'd0; ROM3[1334]<=16'd23832; ROM4[1334]<=16'd57298;
ROM1[1335]<=16'd4819; ROM2[1335]<=16'd0; ROM3[1335]<=16'd23842; ROM4[1335]<=16'd57299;
ROM1[1336]<=16'd4800; ROM2[1336]<=16'd0; ROM3[1336]<=16'd23847; ROM4[1336]<=16'd57293;
ROM1[1337]<=16'd4780; ROM2[1337]<=16'd0; ROM3[1337]<=16'd23843; ROM4[1337]<=16'd57284;
ROM1[1338]<=16'd4765; ROM2[1338]<=16'd0; ROM3[1338]<=16'd23844; ROM4[1338]<=16'd57283;
ROM1[1339]<=16'd4763; ROM2[1339]<=16'd0; ROM3[1339]<=16'd23838; ROM4[1339]<=16'd57286;
ROM1[1340]<=16'd4783; ROM2[1340]<=16'd0; ROM3[1340]<=16'd23832; ROM4[1340]<=16'd57287;
ROM1[1341]<=16'd4838; ROM2[1341]<=16'd0; ROM3[1341]<=16'd23840; ROM4[1341]<=16'd57306;
ROM1[1342]<=16'd4847; ROM2[1342]<=16'd0; ROM3[1342]<=16'd23833; ROM4[1342]<=16'd57307;
ROM1[1343]<=16'd4823; ROM2[1343]<=16'd0; ROM3[1343]<=16'd23831; ROM4[1343]<=16'd57299;
ROM1[1344]<=16'd4799; ROM2[1344]<=16'd0; ROM3[1344]<=16'd23832; ROM4[1344]<=16'd57296;
ROM1[1345]<=16'd4768; ROM2[1345]<=16'd0; ROM3[1345]<=16'd23819; ROM4[1345]<=16'd57276;
ROM1[1346]<=16'd4770; ROM2[1346]<=16'd0; ROM3[1346]<=16'd23838; ROM4[1346]<=16'd57291;
ROM1[1347]<=16'd4769; ROM2[1347]<=16'd0; ROM3[1347]<=16'd23841; ROM4[1347]<=16'd57293;
ROM1[1348]<=16'd4776; ROM2[1348]<=16'd0; ROM3[1348]<=16'd23831; ROM4[1348]<=16'd57285;
ROM1[1349]<=16'd4810; ROM2[1349]<=16'd0; ROM3[1349]<=16'd23825; ROM4[1349]<=16'd57293;
ROM1[1350]<=16'd4845; ROM2[1350]<=16'd0; ROM3[1350]<=16'd23826; ROM4[1350]<=16'd57303;
ROM1[1351]<=16'd4848; ROM2[1351]<=16'd0; ROM3[1351]<=16'd23839; ROM4[1351]<=16'd57313;
ROM1[1352]<=16'd4814; ROM2[1352]<=16'd0; ROM3[1352]<=16'd23826; ROM4[1352]<=16'd57297;
ROM1[1353]<=16'd4790; ROM2[1353]<=16'd0; ROM3[1353]<=16'd23822; ROM4[1353]<=16'd57290;
ROM1[1354]<=16'd4758; ROM2[1354]<=16'd0; ROM3[1354]<=16'd23819; ROM4[1354]<=16'd57282;
ROM1[1355]<=16'd4739; ROM2[1355]<=16'd0; ROM3[1355]<=16'd23812; ROM4[1355]<=16'd57269;
ROM1[1356]<=16'd4748; ROM2[1356]<=16'd0; ROM3[1356]<=16'd23810; ROM4[1356]<=16'd57271;
ROM1[1357]<=16'd4770; ROM2[1357]<=16'd0; ROM3[1357]<=16'd23795; ROM4[1357]<=16'd57266;
ROM1[1358]<=16'd4788; ROM2[1358]<=16'd0; ROM3[1358]<=16'd23770; ROM4[1358]<=16'd57250;
ROM1[1359]<=16'd4784; ROM2[1359]<=16'd0; ROM3[1359]<=16'd23770; ROM4[1359]<=16'd57247;
ROM1[1360]<=16'd4785; ROM2[1360]<=16'd0; ROM3[1360]<=16'd23799; ROM4[1360]<=16'd57268;
ROM1[1361]<=16'd4775; ROM2[1361]<=16'd0; ROM3[1361]<=16'd23814; ROM4[1361]<=16'd57275;
ROM1[1362]<=16'd4752; ROM2[1362]<=16'd0; ROM3[1362]<=16'd23810; ROM4[1362]<=16'd57266;
ROM1[1363]<=16'd4741; ROM2[1363]<=16'd0; ROM3[1363]<=16'd23818; ROM4[1363]<=16'd57271;
ROM1[1364]<=16'd4751; ROM2[1364]<=16'd0; ROM3[1364]<=16'd23827; ROM4[1364]<=16'd57280;
ROM1[1365]<=16'd4785; ROM2[1365]<=16'd0; ROM3[1365]<=16'd23838; ROM4[1365]<=16'd57296;
ROM1[1366]<=16'd4846; ROM2[1366]<=16'd0; ROM3[1366]<=16'd23857; ROM4[1366]<=16'd57324;
ROM1[1367]<=16'd4860; ROM2[1367]<=16'd0; ROM3[1367]<=16'd23860; ROM4[1367]<=16'd57333;
ROM1[1368]<=16'd4808; ROM2[1368]<=16'd0; ROM3[1368]<=16'd23834; ROM4[1368]<=16'd57301;
ROM1[1369]<=16'd4770; ROM2[1369]<=16'd0; ROM3[1369]<=16'd23829; ROM4[1369]<=16'd57284;
ROM1[1370]<=16'd4752; ROM2[1370]<=16'd0; ROM3[1370]<=16'd23832; ROM4[1370]<=16'd57282;
ROM1[1371]<=16'd4750; ROM2[1371]<=16'd0; ROM3[1371]<=16'd23842; ROM4[1371]<=16'd57289;
ROM1[1372]<=16'd4785; ROM2[1372]<=16'd0; ROM3[1372]<=16'd23876; ROM4[1372]<=16'd57322;
ROM1[1373]<=16'd4817; ROM2[1373]<=16'd0; ROM3[1373]<=16'd23887; ROM4[1373]<=16'd57337;
ROM1[1374]<=16'd4825; ROM2[1374]<=16'd0; ROM3[1374]<=16'd23857; ROM4[1374]<=16'd57312;
ROM1[1375]<=16'd4826; ROM2[1375]<=16'd0; ROM3[1375]<=16'd23834; ROM4[1375]<=16'd57297;
ROM1[1376]<=16'd4818; ROM2[1376]<=16'd0; ROM3[1376]<=16'd23831; ROM4[1376]<=16'd57298;
ROM1[1377]<=16'd4801; ROM2[1377]<=16'd0; ROM3[1377]<=16'd23833; ROM4[1377]<=16'd57297;
ROM1[1378]<=16'd4795; ROM2[1378]<=16'd0; ROM3[1378]<=16'd23842; ROM4[1378]<=16'd57306;
ROM1[1379]<=16'd4784; ROM2[1379]<=16'd0; ROM3[1379]<=16'd23852; ROM4[1379]<=16'd57311;
ROM1[1380]<=16'd4779; ROM2[1380]<=16'd0; ROM3[1380]<=16'd23863; ROM4[1380]<=16'd57315;
ROM1[1381]<=16'd4788; ROM2[1381]<=16'd0; ROM3[1381]<=16'd23859; ROM4[1381]<=16'd57313;
ROM1[1382]<=16'd4822; ROM2[1382]<=16'd0; ROM3[1382]<=16'd23858; ROM4[1382]<=16'd57322;
ROM1[1383]<=16'd4860; ROM2[1383]<=16'd0; ROM3[1383]<=16'd23854; ROM4[1383]<=16'd57334;
ROM1[1384]<=16'd4849; ROM2[1384]<=16'd0; ROM3[1384]<=16'd23848; ROM4[1384]<=16'd57327;
ROM1[1385]<=16'd4822; ROM2[1385]<=16'd0; ROM3[1385]<=16'd23851; ROM4[1385]<=16'd57322;
ROM1[1386]<=16'd4804; ROM2[1386]<=16'd0; ROM3[1386]<=16'd23856; ROM4[1386]<=16'd57319;
ROM1[1387]<=16'd4789; ROM2[1387]<=16'd0; ROM3[1387]<=16'd23863; ROM4[1387]<=16'd57315;
ROM1[1388]<=16'd4778; ROM2[1388]<=16'd0; ROM3[1388]<=16'd23869; ROM4[1388]<=16'd57318;
ROM1[1389]<=16'd4776; ROM2[1389]<=16'd0; ROM3[1389]<=16'd23864; ROM4[1389]<=16'd57315;
ROM1[1390]<=16'd4791; ROM2[1390]<=16'd0; ROM3[1390]<=16'd23852; ROM4[1390]<=16'd57309;
ROM1[1391]<=16'd4818; ROM2[1391]<=16'd0; ROM3[1391]<=16'd23838; ROM4[1391]<=16'd57305;
ROM1[1392]<=16'd4829; ROM2[1392]<=16'd0; ROM3[1392]<=16'd23832; ROM4[1392]<=16'd57304;
ROM1[1393]<=16'd4818; ROM2[1393]<=16'd0; ROM3[1393]<=16'd23840; ROM4[1393]<=16'd57307;
ROM1[1394]<=16'd4793; ROM2[1394]<=16'd0; ROM3[1394]<=16'd23846; ROM4[1394]<=16'd57304;
ROM1[1395]<=16'd4775; ROM2[1395]<=16'd0; ROM3[1395]<=16'd23846; ROM4[1395]<=16'd57299;
ROM1[1396]<=16'd4777; ROM2[1396]<=16'd0; ROM3[1396]<=16'd23870; ROM4[1396]<=16'd57318;
ROM1[1397]<=16'd4800; ROM2[1397]<=16'd0; ROM3[1397]<=16'd23894; ROM4[1397]<=16'd57340;
ROM1[1398]<=16'd4811; ROM2[1398]<=16'd0; ROM3[1398]<=16'd23877; ROM4[1398]<=16'd57331;
ROM1[1399]<=16'd4796; ROM2[1399]<=16'd0; ROM3[1399]<=16'd23817; ROM4[1399]<=16'd57281;
ROM1[1400]<=16'd4782; ROM2[1400]<=16'd0; ROM3[1400]<=16'd23774; ROM4[1400]<=16'd57243;
ROM1[1401]<=16'd4762; ROM2[1401]<=16'd0; ROM3[1401]<=16'd23769; ROM4[1401]<=16'd57236;
ROM1[1402]<=16'd4739; ROM2[1402]<=16'd0; ROM3[1402]<=16'd23778; ROM4[1402]<=16'd57238;
ROM1[1403]<=16'd4741; ROM2[1403]<=16'd0; ROM3[1403]<=16'd23806; ROM4[1403]<=16'd57257;
ROM1[1404]<=16'd4734; ROM2[1404]<=16'd0; ROM3[1404]<=16'd23815; ROM4[1404]<=16'd57262;
ROM1[1405]<=16'd4722; ROM2[1405]<=16'd0; ROM3[1405]<=16'd23809; ROM4[1405]<=16'd57257;
ROM1[1406]<=16'd4739; ROM2[1406]<=16'd0; ROM3[1406]<=16'd23813; ROM4[1406]<=16'd57262;
ROM1[1407]<=16'd4778; ROM2[1407]<=16'd0; ROM3[1407]<=16'd23815; ROM4[1407]<=16'd57276;
ROM1[1408]<=16'd4811; ROM2[1408]<=16'd0; ROM3[1408]<=16'd23812; ROM4[1408]<=16'd57283;
ROM1[1409]<=16'd4811; ROM2[1409]<=16'd0; ROM3[1409]<=16'd23814; ROM4[1409]<=16'd57288;
ROM1[1410]<=16'd4804; ROM2[1410]<=16'd0; ROM3[1410]<=16'd23822; ROM4[1410]<=16'd57295;
ROM1[1411]<=16'd4781; ROM2[1411]<=16'd0; ROM3[1411]<=16'd23825; ROM4[1411]<=16'd57292;
ROM1[1412]<=16'd4755; ROM2[1412]<=16'd0; ROM3[1412]<=16'd23820; ROM4[1412]<=16'd57281;
ROM1[1413]<=16'd4748; ROM2[1413]<=16'd0; ROM3[1413]<=16'd23826; ROM4[1413]<=16'd57283;
ROM1[1414]<=16'd4758; ROM2[1414]<=16'd0; ROM3[1414]<=16'd23835; ROM4[1414]<=16'd57291;
ROM1[1415]<=16'd4791; ROM2[1415]<=16'd0; ROM3[1415]<=16'd23838; ROM4[1415]<=16'd57301;
ROM1[1416]<=16'd4830; ROM2[1416]<=16'd0; ROM3[1416]<=16'd23832; ROM4[1416]<=16'd57308;
ROM1[1417]<=16'd4824; ROM2[1417]<=16'd0; ROM3[1417]<=16'd23812; ROM4[1417]<=16'd57290;
ROM1[1418]<=16'd4806; ROM2[1418]<=16'd0; ROM3[1418]<=16'd23816; ROM4[1418]<=16'd57287;
ROM1[1419]<=16'd4809; ROM2[1419]<=16'd0; ROM3[1419]<=16'd23847; ROM4[1419]<=16'd57307;
ROM1[1420]<=16'd4796; ROM2[1420]<=16'd0; ROM3[1420]<=16'd23861; ROM4[1420]<=16'd57313;
ROM1[1421]<=16'd4773; ROM2[1421]<=16'd0; ROM3[1421]<=16'd23863; ROM4[1421]<=16'd57306;
ROM1[1422]<=16'd4753; ROM2[1422]<=16'd0; ROM3[1422]<=16'd23842; ROM4[1422]<=16'd57288;
ROM1[1423]<=16'd4754; ROM2[1423]<=16'd0; ROM3[1423]<=16'd23820; ROM4[1423]<=16'd57273;
ROM1[1424]<=16'd4792; ROM2[1424]<=16'd0; ROM3[1424]<=16'd23815; ROM4[1424]<=16'd57273;
ROM1[1425]<=16'd4812; ROM2[1425]<=16'd0; ROM3[1425]<=16'd23811; ROM4[1425]<=16'd57279;
ROM1[1426]<=16'd4804; ROM2[1426]<=16'd0; ROM3[1426]<=16'd23820; ROM4[1426]<=16'd57285;
ROM1[1427]<=16'd4791; ROM2[1427]<=16'd0; ROM3[1427]<=16'd23832; ROM4[1427]<=16'd57289;
ROM1[1428]<=16'd4784; ROM2[1428]<=16'd0; ROM3[1428]<=16'd23844; ROM4[1428]<=16'd57298;
ROM1[1429]<=16'd4780; ROM2[1429]<=16'd0; ROM3[1429]<=16'd23858; ROM4[1429]<=16'd57306;
ROM1[1430]<=16'd4778; ROM2[1430]<=16'd0; ROM3[1430]<=16'd23867; ROM4[1430]<=16'd57310;
ROM1[1431]<=16'd4784; ROM2[1431]<=16'd0; ROM3[1431]<=16'd23862; ROM4[1431]<=16'd57307;
ROM1[1432]<=16'd4804; ROM2[1432]<=16'd0; ROM3[1432]<=16'd23844; ROM4[1432]<=16'd57303;
ROM1[1433]<=16'd4831; ROM2[1433]<=16'd0; ROM3[1433]<=16'd23834; ROM4[1433]<=16'd57305;
ROM1[1434]<=16'd4831; ROM2[1434]<=16'd0; ROM3[1434]<=16'd23839; ROM4[1434]<=16'd57310;
ROM1[1435]<=16'd4818; ROM2[1435]<=16'd0; ROM3[1435]<=16'd23849; ROM4[1435]<=16'd57316;
ROM1[1436]<=16'd4795; ROM2[1436]<=16'd0; ROM3[1436]<=16'd23853; ROM4[1436]<=16'd57311;
ROM1[1437]<=16'd4771; ROM2[1437]<=16'd0; ROM3[1437]<=16'd23851; ROM4[1437]<=16'd57303;
ROM1[1438]<=16'd4760; ROM2[1438]<=16'd0; ROM3[1438]<=16'd23854; ROM4[1438]<=16'd57304;
ROM1[1439]<=16'd4766; ROM2[1439]<=16'd0; ROM3[1439]<=16'd23859; ROM4[1439]<=16'd57310;
ROM1[1440]<=16'd4788; ROM2[1440]<=16'd0; ROM3[1440]<=16'd23848; ROM4[1440]<=16'd57308;
ROM1[1441]<=16'd4836; ROM2[1441]<=16'd0; ROM3[1441]<=16'd23843; ROM4[1441]<=16'd57315;
ROM1[1442]<=16'd4850; ROM2[1442]<=16'd0; ROM3[1442]<=16'd23850; ROM4[1442]<=16'd57324;
ROM1[1443]<=16'd4820; ROM2[1443]<=16'd0; ROM3[1443]<=16'd23841; ROM4[1443]<=16'd57314;
ROM1[1444]<=16'd4785; ROM2[1444]<=16'd0; ROM3[1444]<=16'd23831; ROM4[1444]<=16'd57296;
ROM1[1445]<=16'd4767; ROM2[1445]<=16'd0; ROM3[1445]<=16'd23834; ROM4[1445]<=16'd57293;
ROM1[1446]<=16'd4745; ROM2[1446]<=16'd0; ROM3[1446]<=16'd23831; ROM4[1446]<=16'd57285;
ROM1[1447]<=16'd4744; ROM2[1447]<=16'd0; ROM3[1447]<=16'd23828; ROM4[1447]<=16'd57282;
ROM1[1448]<=16'd4767; ROM2[1448]<=16'd0; ROM3[1448]<=16'd23830; ROM4[1448]<=16'd57291;
ROM1[1449]<=16'd4788; ROM2[1449]<=16'd0; ROM3[1449]<=16'd23807; ROM4[1449]<=16'd57282;
ROM1[1450]<=16'd4799; ROM2[1450]<=16'd0; ROM3[1450]<=16'd23784; ROM4[1450]<=16'd57267;
ROM1[1451]<=16'd4779; ROM2[1451]<=16'd0; ROM3[1451]<=16'd23774; ROM4[1451]<=16'd57254;
ROM1[1452]<=16'd4756; ROM2[1452]<=16'd0; ROM3[1452]<=16'd23785; ROM4[1452]<=16'd57255;
ROM1[1453]<=16'd4746; ROM2[1453]<=16'd0; ROM3[1453]<=16'd23797; ROM4[1453]<=16'd57260;
ROM1[1454]<=16'd4716; ROM2[1454]<=16'd0; ROM3[1454]<=16'd23791; ROM4[1454]<=16'd57249;
ROM1[1455]<=16'd4706; ROM2[1455]<=16'd0; ROM3[1455]<=16'd23795; ROM4[1455]<=16'd57249;
ROM1[1456]<=16'd4721; ROM2[1456]<=16'd0; ROM3[1456]<=16'd23801; ROM4[1456]<=16'd57258;
ROM1[1457]<=16'd4743; ROM2[1457]<=16'd0; ROM3[1457]<=16'd23791; ROM4[1457]<=16'd57253;
ROM1[1458]<=16'd4773; ROM2[1458]<=16'd0; ROM3[1458]<=16'd23787; ROM4[1458]<=16'd57261;
ROM1[1459]<=16'd4774; ROM2[1459]<=16'd0; ROM3[1459]<=16'd23790; ROM4[1459]<=16'd57266;
ROM1[1460]<=16'd4756; ROM2[1460]<=16'd0; ROM3[1460]<=16'd23799; ROM4[1460]<=16'd57267;
ROM1[1461]<=16'd4742; ROM2[1461]<=16'd0; ROM3[1461]<=16'd23812; ROM4[1461]<=16'd57271;
ROM1[1462]<=16'd4744; ROM2[1462]<=16'd0; ROM3[1462]<=16'd23831; ROM4[1462]<=16'd57281;
ROM1[1463]<=16'd4743; ROM2[1463]<=16'd0; ROM3[1463]<=16'd23848; ROM4[1463]<=16'd57295;
ROM1[1464]<=16'd4765; ROM2[1464]<=16'd0; ROM3[1464]<=16'd23867; ROM4[1464]<=16'd57315;
ROM1[1465]<=16'd4788; ROM2[1465]<=16'd0; ROM3[1465]<=16'd23857; ROM4[1465]<=16'd57311;
ROM1[1466]<=16'd4799; ROM2[1466]<=16'd0; ROM3[1466]<=16'd23827; ROM4[1466]<=16'd57290;
ROM1[1467]<=16'd4822; ROM2[1467]<=16'd0; ROM3[1467]<=16'd23840; ROM4[1467]<=16'd57303;
ROM1[1468]<=16'd4823; ROM2[1468]<=16'd0; ROM3[1468]<=16'd23862; ROM4[1468]<=16'd57319;
ROM1[1469]<=16'd4813; ROM2[1469]<=16'd0; ROM3[1469]<=16'd23878; ROM4[1469]<=16'd57329;
ROM1[1470]<=16'd4798; ROM2[1470]<=16'd0; ROM3[1470]<=16'd23880; ROM4[1470]<=16'd57325;
ROM1[1471]<=16'd4760; ROM2[1471]<=16'd0; ROM3[1471]<=16'd23864; ROM4[1471]<=16'd57301;
ROM1[1472]<=16'd4728; ROM2[1472]<=16'd0; ROM3[1472]<=16'd23836; ROM4[1472]<=16'd57274;
ROM1[1473]<=16'd4735; ROM2[1473]<=16'd0; ROM3[1473]<=16'd23820; ROM4[1473]<=16'd57266;
ROM1[1474]<=16'd4777; ROM2[1474]<=16'd0; ROM3[1474]<=16'd23821; ROM4[1474]<=16'd57275;
ROM1[1475]<=16'd4803; ROM2[1475]<=16'd0; ROM3[1475]<=16'd23820; ROM4[1475]<=16'd57282;
ROM1[1476]<=16'd4802; ROM2[1476]<=16'd0; ROM3[1476]<=16'd23830; ROM4[1476]<=16'd57288;
ROM1[1477]<=16'd4790; ROM2[1477]<=16'd0; ROM3[1477]<=16'd23848; ROM4[1477]<=16'd57297;
ROM1[1478]<=16'd4785; ROM2[1478]<=16'd0; ROM3[1478]<=16'd23866; ROM4[1478]<=16'd57312;
ROM1[1479]<=16'd4769; ROM2[1479]<=16'd0; ROM3[1479]<=16'd23868; ROM4[1479]<=16'd57309;
ROM1[1480]<=16'd4753; ROM2[1480]<=16'd0; ROM3[1480]<=16'd23859; ROM4[1480]<=16'd57299;
ROM1[1481]<=16'd4749; ROM2[1481]<=16'd0; ROM3[1481]<=16'd23846; ROM4[1481]<=16'd57291;
ROM1[1482]<=16'd4768; ROM2[1482]<=16'd0; ROM3[1482]<=16'd23830; ROM4[1482]<=16'd57290;
ROM1[1483]<=16'd4795; ROM2[1483]<=16'd0; ROM3[1483]<=16'd23817; ROM4[1483]<=16'd57288;
ROM1[1484]<=16'd4791; ROM2[1484]<=16'd0; ROM3[1484]<=16'd23816; ROM4[1484]<=16'd57286;
ROM1[1485]<=16'd4777; ROM2[1485]<=16'd0; ROM3[1485]<=16'd23827; ROM4[1485]<=16'd57293;
ROM1[1486]<=16'd4772; ROM2[1486]<=16'd0; ROM3[1486]<=16'd23844; ROM4[1486]<=16'd57304;
ROM1[1487]<=16'd4765; ROM2[1487]<=16'd0; ROM3[1487]<=16'd23859; ROM4[1487]<=16'd57314;
ROM1[1488]<=16'd4748; ROM2[1488]<=16'd0; ROM3[1488]<=16'd23865; ROM4[1488]<=16'd57317;
ROM1[1489]<=16'd4736; ROM2[1489]<=16'd0; ROM3[1489]<=16'd23853; ROM4[1489]<=16'd57299;
ROM1[1490]<=16'd4756; ROM2[1490]<=16'd0; ROM3[1490]<=16'd23845; ROM4[1490]<=16'd57293;
ROM1[1491]<=16'd4802; ROM2[1491]<=16'd0; ROM3[1491]<=16'd23852; ROM4[1491]<=16'd57312;
ROM1[1492]<=16'd4809; ROM2[1492]<=16'd0; ROM3[1492]<=16'd23849; ROM4[1492]<=16'd57313;
ROM1[1493]<=16'd4777; ROM2[1493]<=16'd0; ROM3[1493]<=16'd23833; ROM4[1493]<=16'd57294;
ROM1[1494]<=16'd4751; ROM2[1494]<=16'd0; ROM3[1494]<=16'd23829; ROM4[1494]<=16'd57287;
ROM1[1495]<=16'd4740; ROM2[1495]<=16'd0; ROM3[1495]<=16'd23834; ROM4[1495]<=16'd57285;
ROM1[1496]<=16'd4730; ROM2[1496]<=16'd0; ROM3[1496]<=16'd23841; ROM4[1496]<=16'd57286;
ROM1[1497]<=16'd4725; ROM2[1497]<=16'd0; ROM3[1497]<=16'd23840; ROM4[1497]<=16'd57286;
ROM1[1498]<=16'd4731; ROM2[1498]<=16'd0; ROM3[1498]<=16'd23829; ROM4[1498]<=16'd57276;
ROM1[1499]<=16'd4753; ROM2[1499]<=16'd0; ROM3[1499]<=16'd23807; ROM4[1499]<=16'd57266;
ROM1[1500]<=16'd4770; ROM2[1500]<=16'd0; ROM3[1500]<=16'd23796; ROM4[1500]<=16'd57262;
ROM1[1501]<=16'd4775; ROM2[1501]<=16'd0; ROM3[1501]<=16'd23809; ROM4[1501]<=16'd57274;
ROM1[1502]<=16'd4764; ROM2[1502]<=16'd0; ROM3[1502]<=16'd23819; ROM4[1502]<=16'd57282;
ROM1[1503]<=16'd4747; ROM2[1503]<=16'd0; ROM3[1503]<=16'd23825; ROM4[1503]<=16'd57283;
ROM1[1504]<=16'd4738; ROM2[1504]<=16'd0; ROM3[1504]<=16'd23835; ROM4[1504]<=16'd57290;
ROM1[1505]<=16'd4739; ROM2[1505]<=16'd0; ROM3[1505]<=16'd23843; ROM4[1505]<=16'd57295;
ROM1[1506]<=16'd4739; ROM2[1506]<=16'd0; ROM3[1506]<=16'd23831; ROM4[1506]<=16'd57281;
ROM1[1507]<=16'd4754; ROM2[1507]<=16'd0; ROM3[1507]<=16'd23805; ROM4[1507]<=16'd57264;
ROM1[1508]<=16'd4777; ROM2[1508]<=16'd0; ROM3[1508]<=16'd23794; ROM4[1508]<=16'd57259;
ROM1[1509]<=16'd4771; ROM2[1509]<=16'd0; ROM3[1509]<=16'd23798; ROM4[1509]<=16'd57263;
ROM1[1510]<=16'd4757; ROM2[1510]<=16'd0; ROM3[1510]<=16'd23810; ROM4[1510]<=16'd57269;
ROM1[1511]<=16'd4753; ROM2[1511]<=16'd0; ROM3[1511]<=16'd23832; ROM4[1511]<=16'd57282;
ROM1[1512]<=16'd4769; ROM2[1512]<=16'd0; ROM3[1512]<=16'd23863; ROM4[1512]<=16'd57307;
ROM1[1513]<=16'd4782; ROM2[1513]<=16'd0; ROM3[1513]<=16'd23892; ROM4[1513]<=16'd57328;
ROM1[1514]<=16'd4769; ROM2[1514]<=16'd0; ROM3[1514]<=16'd23878; ROM4[1514]<=16'd57315;
ROM1[1515]<=16'd4758; ROM2[1515]<=16'd0; ROM3[1515]<=16'd23834; ROM4[1515]<=16'd57280;
ROM1[1516]<=16'd4775; ROM2[1516]<=16'd0; ROM3[1516]<=16'd23807; ROM4[1516]<=16'd57265;
ROM1[1517]<=16'd4766; ROM2[1517]<=16'd0; ROM3[1517]<=16'd23782; ROM4[1517]<=16'd57253;
ROM1[1518]<=16'd4758; ROM2[1518]<=16'd0; ROM3[1518]<=16'd23792; ROM4[1518]<=16'd57258;
ROM1[1519]<=16'd4760; ROM2[1519]<=16'd0; ROM3[1519]<=16'd23829; ROM4[1519]<=16'd57286;
ROM1[1520]<=16'd4735; ROM2[1520]<=16'd0; ROM3[1520]<=16'd23824; ROM4[1520]<=16'd57280;
ROM1[1521]<=16'd4701; ROM2[1521]<=16'd0; ROM3[1521]<=16'd23809; ROM4[1521]<=16'd57258;
ROM1[1522]<=16'd4695; ROM2[1522]<=16'd0; ROM3[1522]<=16'd23811; ROM4[1522]<=16'd57258;
ROM1[1523]<=16'd4704; ROM2[1523]<=16'd0; ROM3[1523]<=16'd23790; ROM4[1523]<=16'd57246;
ROM1[1524]<=16'd4720; ROM2[1524]<=16'd0; ROM3[1524]<=16'd23758; ROM4[1524]<=16'd57225;
ROM1[1525]<=16'd4743; ROM2[1525]<=16'd0; ROM3[1525]<=16'd23755; ROM4[1525]<=16'd57230;
ROM1[1526]<=16'd4755; ROM2[1526]<=16'd0; ROM3[1526]<=16'd23779; ROM4[1526]<=16'd57254;
ROM1[1527]<=16'd4767; ROM2[1527]<=16'd0; ROM3[1527]<=16'd23817; ROM4[1527]<=16'd57281;
ROM1[1528]<=16'd4786; ROM2[1528]<=16'd0; ROM3[1528]<=16'd23853; ROM4[1528]<=16'd57311;
ROM1[1529]<=16'd4782; ROM2[1529]<=16'd0; ROM3[1529]<=16'd23866; ROM4[1529]<=16'd57321;
ROM1[1530]<=16'd4765; ROM2[1530]<=16'd0; ROM3[1530]<=16'd23863; ROM4[1530]<=16'd57312;
ROM1[1531]<=16'd4765; ROM2[1531]<=16'd0; ROM3[1531]<=16'd23859; ROM4[1531]<=16'd57312;
ROM1[1532]<=16'd4803; ROM2[1532]<=16'd0; ROM3[1532]<=16'd23870; ROM4[1532]<=16'd57326;
ROM1[1533]<=16'd4845; ROM2[1533]<=16'd0; ROM3[1533]<=16'd23878; ROM4[1533]<=16'd57336;
ROM1[1534]<=16'd4827; ROM2[1534]<=16'd0; ROM3[1534]<=16'd23861; ROM4[1534]<=16'd57319;
ROM1[1535]<=16'd4799; ROM2[1535]<=16'd0; ROM3[1535]<=16'd23854; ROM4[1535]<=16'd57305;
ROM1[1536]<=16'd4780; ROM2[1536]<=16'd0; ROM3[1536]<=16'd23863; ROM4[1536]<=16'd57305;
ROM1[1537]<=16'd4765; ROM2[1537]<=16'd0; ROM3[1537]<=16'd23869; ROM4[1537]<=16'd57307;
ROM1[1538]<=16'd4749; ROM2[1538]<=16'd0; ROM3[1538]<=16'd23874; ROM4[1538]<=16'd57312;
ROM1[1539]<=16'd4753; ROM2[1539]<=16'd0; ROM3[1539]<=16'd23879; ROM4[1539]<=16'd57316;
ROM1[1540]<=16'd4774; ROM2[1540]<=16'd0; ROM3[1540]<=16'd23870; ROM4[1540]<=16'd57315;
ROM1[1541]<=16'd4801; ROM2[1541]<=16'd0; ROM3[1541]<=16'd23847; ROM4[1541]<=16'd57308;
ROM1[1542]<=16'd4811; ROM2[1542]<=16'd0; ROM3[1542]<=16'd23840; ROM4[1542]<=16'd57306;
ROM1[1543]<=16'd4794; ROM2[1543]<=16'd0; ROM3[1543]<=16'd23841; ROM4[1543]<=16'd57307;
ROM1[1544]<=16'd4758; ROM2[1544]<=16'd0; ROM3[1544]<=16'd23834; ROM4[1544]<=16'd57297;
ROM1[1545]<=16'd4744; ROM2[1545]<=16'd0; ROM3[1545]<=16'd23842; ROM4[1545]<=16'd57297;
ROM1[1546]<=16'd4744; ROM2[1546]<=16'd0; ROM3[1546]<=16'd23859; ROM4[1546]<=16'd57306;
ROM1[1547]<=16'd4747; ROM2[1547]<=16'd0; ROM3[1547]<=16'd23862; ROM4[1547]<=16'd57306;
ROM1[1548]<=16'd4756; ROM2[1548]<=16'd0; ROM3[1548]<=16'd23843; ROM4[1548]<=16'd57298;
ROM1[1549]<=16'd4804; ROM2[1549]<=16'd0; ROM3[1549]<=16'd23846; ROM4[1549]<=16'd57315;
ROM1[1550]<=16'd4857; ROM2[1550]<=16'd0; ROM3[1550]<=16'd23873; ROM4[1550]<=16'd57347;
ROM1[1551]<=16'd4830; ROM2[1551]<=16'd0; ROM3[1551]<=16'd23861; ROM4[1551]<=16'd57330;
ROM1[1552]<=16'd4779; ROM2[1552]<=16'd0; ROM3[1552]<=16'd23833; ROM4[1552]<=16'd57292;
ROM1[1553]<=16'd4759; ROM2[1553]<=16'd0; ROM3[1553]<=16'd23834; ROM4[1553]<=16'd57285;
ROM1[1554]<=16'd4736; ROM2[1554]<=16'd0; ROM3[1554]<=16'd23833; ROM4[1554]<=16'd57282;
ROM1[1555]<=16'd4724; ROM2[1555]<=16'd0; ROM3[1555]<=16'd23832; ROM4[1555]<=16'd57276;
ROM1[1556]<=16'd4742; ROM2[1556]<=16'd0; ROM3[1556]<=16'd23836; ROM4[1556]<=16'd57281;
ROM1[1557]<=16'd4751; ROM2[1557]<=16'd0; ROM3[1557]<=16'd23812; ROM4[1557]<=16'd57269;
ROM1[1558]<=16'd4765; ROM2[1558]<=16'd0; ROM3[1558]<=16'd23787; ROM4[1558]<=16'd57253;
ROM1[1559]<=16'd4778; ROM2[1559]<=16'd0; ROM3[1559]<=16'd23800; ROM4[1559]<=16'd57266;
ROM1[1560]<=16'd4786; ROM2[1560]<=16'd0; ROM3[1560]<=16'd23831; ROM4[1560]<=16'd57293;
ROM1[1561]<=16'd4784; ROM2[1561]<=16'd0; ROM3[1561]<=16'd23850; ROM4[1561]<=16'd57308;
ROM1[1562]<=16'd4760; ROM2[1562]<=16'd0; ROM3[1562]<=16'd23844; ROM4[1562]<=16'd57299;
ROM1[1563]<=16'd4738; ROM2[1563]<=16'd0; ROM3[1563]<=16'd23839; ROM4[1563]<=16'd57289;
ROM1[1564]<=16'd4721; ROM2[1564]<=16'd0; ROM3[1564]<=16'd23820; ROM4[1564]<=16'd57270;
ROM1[1565]<=16'd4730; ROM2[1565]<=16'd0; ROM3[1565]<=16'd23797; ROM4[1565]<=16'd57258;
ROM1[1566]<=16'd4782; ROM2[1566]<=16'd0; ROM3[1566]<=16'd23804; ROM4[1566]<=16'd57274;
ROM1[1567]<=16'd4812; ROM2[1567]<=16'd0; ROM3[1567]<=16'd23823; ROM4[1567]<=16'd57296;
ROM1[1568]<=16'd4790; ROM2[1568]<=16'd0; ROM3[1568]<=16'd23825; ROM4[1568]<=16'd57293;
ROM1[1569]<=16'd4764; ROM2[1569]<=16'd0; ROM3[1569]<=16'd23826; ROM4[1569]<=16'd57285;
ROM1[1570]<=16'd4767; ROM2[1570]<=16'd0; ROM3[1570]<=16'd23840; ROM4[1570]<=16'd57294;
ROM1[1571]<=16'd4748; ROM2[1571]<=16'd0; ROM3[1571]<=16'd23841; ROM4[1571]<=16'd57288;
ROM1[1572]<=16'd4733; ROM2[1572]<=16'd0; ROM3[1572]<=16'd23827; ROM4[1572]<=16'd57275;
ROM1[1573]<=16'd4759; ROM2[1573]<=16'd0; ROM3[1573]<=16'd23830; ROM4[1573]<=16'd57284;
ROM1[1574]<=16'd4777; ROM2[1574]<=16'd0; ROM3[1574]<=16'd23811; ROM4[1574]<=16'd57275;
ROM1[1575]<=16'd4762; ROM2[1575]<=16'd0; ROM3[1575]<=16'd23778; ROM4[1575]<=16'd57248;
ROM1[1576]<=16'd4766; ROM2[1576]<=16'd0; ROM3[1576]<=16'd23798; ROM4[1576]<=16'd57262;
ROM1[1577]<=16'd4768; ROM2[1577]<=16'd0; ROM3[1577]<=16'd23830; ROM4[1577]<=16'd57285;
ROM1[1578]<=16'd4762; ROM2[1578]<=16'd0; ROM3[1578]<=16'd23846; ROM4[1578]<=16'd57300;
ROM1[1579]<=16'd4760; ROM2[1579]<=16'd0; ROM3[1579]<=16'd23865; ROM4[1579]<=16'd57314;
ROM1[1580]<=16'd4754; ROM2[1580]<=16'd0; ROM3[1580]<=16'd23874; ROM4[1580]<=16'd57314;
ROM1[1581]<=16'd4764; ROM2[1581]<=16'd0; ROM3[1581]<=16'd23873; ROM4[1581]<=16'd57315;
ROM1[1582]<=16'd4790; ROM2[1582]<=16'd0; ROM3[1582]<=16'd23864; ROM4[1582]<=16'd57316;
ROM1[1583]<=16'd4799; ROM2[1583]<=16'd0; ROM3[1583]<=16'd23837; ROM4[1583]<=16'd57301;
ROM1[1584]<=16'd4795; ROM2[1584]<=16'd0; ROM3[1584]<=16'd23836; ROM4[1584]<=16'd57302;
ROM1[1585]<=16'd4777; ROM2[1585]<=16'd0; ROM3[1585]<=16'd23845; ROM4[1585]<=16'd57299;
ROM1[1586]<=16'd4761; ROM2[1586]<=16'd0; ROM3[1586]<=16'd23856; ROM4[1586]<=16'd57302;
ROM1[1587]<=16'd4787; ROM2[1587]<=16'd0; ROM3[1587]<=16'd23904; ROM4[1587]<=16'd57343;
ROM1[1588]<=16'd4785; ROM2[1588]<=16'd0; ROM3[1588]<=16'd23916; ROM4[1588]<=16'd57350;
ROM1[1589]<=16'd4758; ROM2[1589]<=16'd0; ROM3[1589]<=16'd23879; ROM4[1589]<=16'd57319;
ROM1[1590]<=16'd4764; ROM2[1590]<=16'd0; ROM3[1590]<=16'd23849; ROM4[1590]<=16'd57296;
ROM1[1591]<=16'd4796; ROM2[1591]<=16'd0; ROM3[1591]<=16'd23836; ROM4[1591]<=16'd57298;
ROM1[1592]<=16'd4814; ROM2[1592]<=16'd0; ROM3[1592]<=16'd23839; ROM4[1592]<=16'd57307;
ROM1[1593]<=16'd4799; ROM2[1593]<=16'd0; ROM3[1593]<=16'd23846; ROM4[1593]<=16'd57307;
ROM1[1594]<=16'd4782; ROM2[1594]<=16'd0; ROM3[1594]<=16'd23860; ROM4[1594]<=16'd57309;
ROM1[1595]<=16'd4768; ROM2[1595]<=16'd0; ROM3[1595]<=16'd23858; ROM4[1595]<=16'd57304;
ROM1[1596]<=16'd4748; ROM2[1596]<=16'd0; ROM3[1596]<=16'd23859; ROM4[1596]<=16'd57303;
ROM1[1597]<=16'd4748; ROM2[1597]<=16'd0; ROM3[1597]<=16'd23867; ROM4[1597]<=16'd57307;
ROM1[1598]<=16'd4765; ROM2[1598]<=16'd0; ROM3[1598]<=16'd23862; ROM4[1598]<=16'd57309;
ROM1[1599]<=16'd4792; ROM2[1599]<=16'd0; ROM3[1599]<=16'd23844; ROM4[1599]<=16'd57301;
ROM1[1600]<=16'd4807; ROM2[1600]<=16'd0; ROM3[1600]<=16'd23830; ROM4[1600]<=16'd57291;
ROM1[1601]<=16'd4797; ROM2[1601]<=16'd0; ROM3[1601]<=16'd23831; ROM4[1601]<=16'd57290;
ROM1[1602]<=16'd4785; ROM2[1602]<=16'd0; ROM3[1602]<=16'd23844; ROM4[1602]<=16'd57297;
ROM1[1603]<=16'd4788; ROM2[1603]<=16'd0; ROM3[1603]<=16'd23869; ROM4[1603]<=16'd57315;
ROM1[1604]<=16'd4772; ROM2[1604]<=16'd0; ROM3[1604]<=16'd23875; ROM4[1604]<=16'd57317;
ROM1[1605]<=16'd4733; ROM2[1605]<=16'd0; ROM3[1605]<=16'd23845; ROM4[1605]<=16'd57285;
ROM1[1606]<=16'd4728; ROM2[1606]<=16'd0; ROM3[1606]<=16'd23826; ROM4[1606]<=16'd57265;
ROM1[1607]<=16'd4749; ROM2[1607]<=16'd0; ROM3[1607]<=16'd23807; ROM4[1607]<=16'd57260;
ROM1[1608]<=16'd4786; ROM2[1608]<=16'd0; ROM3[1608]<=16'd23807; ROM4[1608]<=16'd57269;
ROM1[1609]<=16'd4826; ROM2[1609]<=16'd0; ROM3[1609]<=16'd23849; ROM4[1609]<=16'd57308;
ROM1[1610]<=16'd4803; ROM2[1610]<=16'd0; ROM3[1610]<=16'd23850; ROM4[1610]<=16'd57305;
ROM1[1611]<=16'd4756; ROM2[1611]<=16'd0; ROM3[1611]<=16'd23822; ROM4[1611]<=16'd57268;
ROM1[1612]<=16'd4736; ROM2[1612]<=16'd0; ROM3[1612]<=16'd23815; ROM4[1612]<=16'd57257;
ROM1[1613]<=16'd4717; ROM2[1613]<=16'd0; ROM3[1613]<=16'd23809; ROM4[1613]<=16'd57253;
ROM1[1614]<=16'd4723; ROM2[1614]<=16'd0; ROM3[1614]<=16'd23806; ROM4[1614]<=16'd57254;
ROM1[1615]<=16'd4747; ROM2[1615]<=16'd0; ROM3[1615]<=16'd23808; ROM4[1615]<=16'd57257;
ROM1[1616]<=16'd4772; ROM2[1616]<=16'd0; ROM3[1616]<=16'd23796; ROM4[1616]<=16'd57256;
ROM1[1617]<=16'd4783; ROM2[1617]<=16'd0; ROM3[1617]<=16'd23791; ROM4[1617]<=16'd57258;
ROM1[1618]<=16'd4763; ROM2[1618]<=16'd0; ROM3[1618]<=16'd23786; ROM4[1618]<=16'd57253;
ROM1[1619]<=16'd4765; ROM2[1619]<=16'd0; ROM3[1619]<=16'd23814; ROM4[1619]<=16'd57273;
ROM1[1620]<=16'd4764; ROM2[1620]<=16'd0; ROM3[1620]<=16'd23832; ROM4[1620]<=16'd57281;
ROM1[1621]<=16'd4725; ROM2[1621]<=16'd0; ROM3[1621]<=16'd23817; ROM4[1621]<=16'd57254;
ROM1[1622]<=16'd4712; ROM2[1622]<=16'd0; ROM3[1622]<=16'd23816; ROM4[1622]<=16'd57243;
ROM1[1623]<=16'd4714; ROM2[1623]<=16'd0; ROM3[1623]<=16'd23798; ROM4[1623]<=16'd57233;
ROM1[1624]<=16'd4740; ROM2[1624]<=16'd0; ROM3[1624]<=16'd23782; ROM4[1624]<=16'd57225;
ROM1[1625]<=16'd4768; ROM2[1625]<=16'd0; ROM3[1625]<=16'd23783; ROM4[1625]<=16'd57236;
ROM1[1626]<=16'd4761; ROM2[1626]<=16'd0; ROM3[1626]<=16'd23796; ROM4[1626]<=16'd57245;
ROM1[1627]<=16'd4742; ROM2[1627]<=16'd0; ROM3[1627]<=16'd23805; ROM4[1627]<=16'd57247;
ROM1[1628]<=16'd4735; ROM2[1628]<=16'd0; ROM3[1628]<=16'd23818; ROM4[1628]<=16'd57259;
ROM1[1629]<=16'd4723; ROM2[1629]<=16'd0; ROM3[1629]<=16'd23832; ROM4[1629]<=16'd57264;
ROM1[1630]<=16'd4724; ROM2[1630]<=16'd0; ROM3[1630]<=16'd23838; ROM4[1630]<=16'd57270;
ROM1[1631]<=16'd4752; ROM2[1631]<=16'd0; ROM3[1631]<=16'd23848; ROM4[1631]<=16'd57285;
ROM1[1632]<=16'd4777; ROM2[1632]<=16'd0; ROM3[1632]<=16'd23835; ROM4[1632]<=16'd57284;
ROM1[1633]<=16'd4798; ROM2[1633]<=16'd0; ROM3[1633]<=16'd23821; ROM4[1633]<=16'd57284;
ROM1[1634]<=16'd4796; ROM2[1634]<=16'd0; ROM3[1634]<=16'd23823; ROM4[1634]<=16'd57284;
ROM1[1635]<=16'd4781; ROM2[1635]<=16'd0; ROM3[1635]<=16'd23830; ROM4[1635]<=16'd57283;
ROM1[1636]<=16'd4777; ROM2[1636]<=16'd0; ROM3[1636]<=16'd23852; ROM4[1636]<=16'd57301;
ROM1[1637]<=16'd4781; ROM2[1637]<=16'd0; ROM3[1637]<=16'd23872; ROM4[1637]<=16'd57318;
ROM1[1638]<=16'd4768; ROM2[1638]<=16'd0; ROM3[1638]<=16'd23874; ROM4[1638]<=16'd57316;
ROM1[1639]<=16'd4761; ROM2[1639]<=16'd0; ROM3[1639]<=16'd23863; ROM4[1639]<=16'd57304;
ROM1[1640]<=16'd4777; ROM2[1640]<=16'd0; ROM3[1640]<=16'd23846; ROM4[1640]<=16'd57291;
ROM1[1641]<=16'd4813; ROM2[1641]<=16'd0; ROM3[1641]<=16'd23836; ROM4[1641]<=16'd57293;
ROM1[1642]<=16'd4839; ROM2[1642]<=16'd0; ROM3[1642]<=16'd23846; ROM4[1642]<=16'd57311;
ROM1[1643]<=16'd4825; ROM2[1643]<=16'd0; ROM3[1643]<=16'd23851; ROM4[1643]<=16'd57312;
ROM1[1644]<=16'd4796; ROM2[1644]<=16'd0; ROM3[1644]<=16'd23855; ROM4[1644]<=16'd57305;
ROM1[1645]<=16'd4773; ROM2[1645]<=16'd0; ROM3[1645]<=16'd23859; ROM4[1645]<=16'd57302;
ROM1[1646]<=16'd4756; ROM2[1646]<=16'd0; ROM3[1646]<=16'd23859; ROM4[1646]<=16'd57299;
ROM1[1647]<=16'd4766; ROM2[1647]<=16'd0; ROM3[1647]<=16'd23864; ROM4[1647]<=16'd57304;
ROM1[1648]<=16'd4788; ROM2[1648]<=16'd0; ROM3[1648]<=16'd23857; ROM4[1648]<=16'd57304;
ROM1[1649]<=16'd4833; ROM2[1649]<=16'd0; ROM3[1649]<=16'd23850; ROM4[1649]<=16'd57316;
ROM1[1650]<=16'd4871; ROM2[1650]<=16'd0; ROM3[1650]<=16'd23860; ROM4[1650]<=16'd57335;
ROM1[1651]<=16'd4859; ROM2[1651]<=16'd0; ROM3[1651]<=16'd23867; ROM4[1651]<=16'd57339;
ROM1[1652]<=16'd4829; ROM2[1652]<=16'd0; ROM3[1652]<=16'd23862; ROM4[1652]<=16'd57331;
ROM1[1653]<=16'd4811; ROM2[1653]<=16'd0; ROM3[1653]<=16'd23866; ROM4[1653]<=16'd57329;
ROM1[1654]<=16'd4778; ROM2[1654]<=16'd0; ROM3[1654]<=16'd23855; ROM4[1654]<=16'd57312;
ROM1[1655]<=16'd4749; ROM2[1655]<=16'd0; ROM3[1655]<=16'd23835; ROM4[1655]<=16'd57289;
ROM1[1656]<=16'd4772; ROM2[1656]<=16'd0; ROM3[1656]<=16'd23841; ROM4[1656]<=16'd57296;
ROM1[1657]<=16'd4803; ROM2[1657]<=16'd0; ROM3[1657]<=16'd23833; ROM4[1657]<=16'd57295;
ROM1[1658]<=16'd4822; ROM2[1658]<=16'd0; ROM3[1658]<=16'd23814; ROM4[1658]<=16'd57285;
ROM1[1659]<=16'd4822; ROM2[1659]<=16'd0; ROM3[1659]<=16'd23818; ROM4[1659]<=16'd57291;
ROM1[1660]<=16'd4811; ROM2[1660]<=16'd0; ROM3[1660]<=16'd23830; ROM4[1660]<=16'd57299;
ROM1[1661]<=16'd4793; ROM2[1661]<=16'd0; ROM3[1661]<=16'd23839; ROM4[1661]<=16'd57298;
ROM1[1662]<=16'd4769; ROM2[1662]<=16'd0; ROM3[1662]<=16'd23835; ROM4[1662]<=16'd57290;
ROM1[1663]<=16'd4751; ROM2[1663]<=16'd0; ROM3[1663]<=16'd23840; ROM4[1663]<=16'd57290;
ROM1[1664]<=16'd4754; ROM2[1664]<=16'd0; ROM3[1664]<=16'd23845; ROM4[1664]<=16'd57298;
ROM1[1665]<=16'd4776; ROM2[1665]<=16'd0; ROM3[1665]<=16'd23838; ROM4[1665]<=16'd57301;
ROM1[1666]<=16'd4809; ROM2[1666]<=16'd0; ROM3[1666]<=16'd23827; ROM4[1666]<=16'd57300;
ROM1[1667]<=16'd4818; ROM2[1667]<=16'd0; ROM3[1667]<=16'd23820; ROM4[1667]<=16'd57301;
ROM1[1668]<=16'd4788; ROM2[1668]<=16'd0; ROM3[1668]<=16'd23811; ROM4[1668]<=16'd57285;
ROM1[1669]<=16'd4761; ROM2[1669]<=16'd0; ROM3[1669]<=16'd23807; ROM4[1669]<=16'd57276;
ROM1[1670]<=16'd4753; ROM2[1670]<=16'd0; ROM3[1670]<=16'd23821; ROM4[1670]<=16'd57284;
ROM1[1671]<=16'd4737; ROM2[1671]<=16'd0; ROM3[1671]<=16'd23829; ROM4[1671]<=16'd57282;
ROM1[1672]<=16'd4730; ROM2[1672]<=16'd0; ROM3[1672]<=16'd23823; ROM4[1672]<=16'd57274;
ROM1[1673]<=16'd4753; ROM2[1673]<=16'd0; ROM3[1673]<=16'd23822; ROM4[1673]<=16'd57277;
ROM1[1674]<=16'd4787; ROM2[1674]<=16'd0; ROM3[1674]<=16'd23811; ROM4[1674]<=16'd57277;
ROM1[1675]<=16'd4797; ROM2[1675]<=16'd0; ROM3[1675]<=16'd23796; ROM4[1675]<=16'd57271;
ROM1[1676]<=16'd4776; ROM2[1676]<=16'd0; ROM3[1676]<=16'd23788; ROM4[1676]<=16'd57259;
ROM1[1677]<=16'd4748; ROM2[1677]<=16'd0; ROM3[1677]<=16'd23785; ROM4[1677]<=16'd57248;
ROM1[1678]<=16'd4729; ROM2[1678]<=16'd0; ROM3[1678]<=16'd23786; ROM4[1678]<=16'd57242;
ROM1[1679]<=16'd4722; ROM2[1679]<=16'd0; ROM3[1679]<=16'd23796; ROM4[1679]<=16'd57244;
ROM1[1680]<=16'd4724; ROM2[1680]<=16'd0; ROM3[1680]<=16'd23805; ROM4[1680]<=16'd57255;
ROM1[1681]<=16'd4732; ROM2[1681]<=16'd0; ROM3[1681]<=16'd23800; ROM4[1681]<=16'd57258;
ROM1[1682]<=16'd4757; ROM2[1682]<=16'd0; ROM3[1682]<=16'd23786; ROM4[1682]<=16'd57253;
ROM1[1683]<=16'd4777; ROM2[1683]<=16'd0; ROM3[1683]<=16'd23767; ROM4[1683]<=16'd57247;
ROM1[1684]<=16'd4775; ROM2[1684]<=16'd0; ROM3[1684]<=16'd23769; ROM4[1684]<=16'd57245;
ROM1[1685]<=16'd4757; ROM2[1685]<=16'd0; ROM3[1685]<=16'd23776; ROM4[1685]<=16'd57242;
ROM1[1686]<=16'd4738; ROM2[1686]<=16'd0; ROM3[1686]<=16'd23785; ROM4[1686]<=16'd57243;
ROM1[1687]<=16'd4724; ROM2[1687]<=16'd0; ROM3[1687]<=16'd23789; ROM4[1687]<=16'd57245;
ROM1[1688]<=16'd4723; ROM2[1688]<=16'd0; ROM3[1688]<=16'd23798; ROM4[1688]<=16'd57252;
ROM1[1689]<=16'd4751; ROM2[1689]<=16'd0; ROM3[1689]<=16'd23815; ROM4[1689]<=16'd57270;
ROM1[1690]<=16'd4783; ROM2[1690]<=16'd0; ROM3[1690]<=16'd23817; ROM4[1690]<=16'd57279;
ROM1[1691]<=16'd4805; ROM2[1691]<=16'd0; ROM3[1691]<=16'd23801; ROM4[1691]<=16'd57275;
ROM1[1692]<=16'd4796; ROM2[1692]<=16'd0; ROM3[1692]<=16'd23787; ROM4[1692]<=16'd57262;
ROM1[1693]<=16'd4770; ROM2[1693]<=16'd0; ROM3[1693]<=16'd23782; ROM4[1693]<=16'd57252;
ROM1[1694]<=16'd4743; ROM2[1694]<=16'd0; ROM3[1694]<=16'd23781; ROM4[1694]<=16'd57244;
ROM1[1695]<=16'd4735; ROM2[1695]<=16'd0; ROM3[1695]<=16'd23789; ROM4[1695]<=16'd57245;
ROM1[1696]<=16'd4733; ROM2[1696]<=16'd0; ROM3[1696]<=16'd23810; ROM4[1696]<=16'd57261;
ROM1[1697]<=16'd4747; ROM2[1697]<=16'd0; ROM3[1697]<=16'd23828; ROM4[1697]<=16'd57280;
ROM1[1698]<=16'd4768; ROM2[1698]<=16'd0; ROM3[1698]<=16'd23826; ROM4[1698]<=16'd57284;
ROM1[1699]<=16'd4802; ROM2[1699]<=16'd0; ROM3[1699]<=16'd23818; ROM4[1699]<=16'd57287;
ROM1[1700]<=16'd4807; ROM2[1700]<=16'd0; ROM3[1700]<=16'd23800; ROM4[1700]<=16'd57276;
ROM1[1701]<=16'd4766; ROM2[1701]<=16'd0; ROM3[1701]<=16'd23778; ROM4[1701]<=16'd57249;
ROM1[1702]<=16'd4751; ROM2[1702]<=16'd0; ROM3[1702]<=16'd23787; ROM4[1702]<=16'd57252;
ROM1[1703]<=16'd4757; ROM2[1703]<=16'd0; ROM3[1703]<=16'd23813; ROM4[1703]<=16'd57270;
ROM1[1704]<=16'd4757; ROM2[1704]<=16'd0; ROM3[1704]<=16'd23832; ROM4[1704]<=16'd57282;
ROM1[1705]<=16'd4750; ROM2[1705]<=16'd0; ROM3[1705]<=16'd23837; ROM4[1705]<=16'd57285;
ROM1[1706]<=16'd4754; ROM2[1706]<=16'd0; ROM3[1706]<=16'd23838; ROM4[1706]<=16'd57283;
ROM1[1707]<=16'd4787; ROM2[1707]<=16'd0; ROM3[1707]<=16'd23829; ROM4[1707]<=16'd57287;
ROM1[1708]<=16'd4813; ROM2[1708]<=16'd0; ROM3[1708]<=16'd23812; ROM4[1708]<=16'd57285;
ROM1[1709]<=16'd4807; ROM2[1709]<=16'd0; ROM3[1709]<=16'd23813; ROM4[1709]<=16'd57286;
ROM1[1710]<=16'd4794; ROM2[1710]<=16'd0; ROM3[1710]<=16'd23825; ROM4[1710]<=16'd57293;
ROM1[1711]<=16'd4783; ROM2[1711]<=16'd0; ROM3[1711]<=16'd23838; ROM4[1711]<=16'd57298;
ROM1[1712]<=16'd4775; ROM2[1712]<=16'd0; ROM3[1712]<=16'd23855; ROM4[1712]<=16'd57307;
ROM1[1713]<=16'd4751; ROM2[1713]<=16'd0; ROM3[1713]<=16'd23847; ROM4[1713]<=16'd57291;
ROM1[1714]<=16'd4754; ROM2[1714]<=16'd0; ROM3[1714]<=16'd23838; ROM4[1714]<=16'd57285;
ROM1[1715]<=16'd4780; ROM2[1715]<=16'd0; ROM3[1715]<=16'd23833; ROM4[1715]<=16'd57288;
ROM1[1716]<=16'd4813; ROM2[1716]<=16'd0; ROM3[1716]<=16'd23824; ROM4[1716]<=16'd57287;
ROM1[1717]<=16'd4825; ROM2[1717]<=16'd0; ROM3[1717]<=16'd23823; ROM4[1717]<=16'd57293;
ROM1[1718]<=16'd4800; ROM2[1718]<=16'd0; ROM3[1718]<=16'd23825; ROM4[1718]<=16'd57290;
ROM1[1719]<=16'd4779; ROM2[1719]<=16'd0; ROM3[1719]<=16'd23831; ROM4[1719]<=16'd57289;
ROM1[1720]<=16'd4773; ROM2[1720]<=16'd0; ROM3[1720]<=16'd23837; ROM4[1720]<=16'd57293;
ROM1[1721]<=16'd4765; ROM2[1721]<=16'd0; ROM3[1721]<=16'd23850; ROM4[1721]<=16'd57300;
ROM1[1722]<=16'd4772; ROM2[1722]<=16'd0; ROM3[1722]<=16'd23856; ROM4[1722]<=16'd57306;
ROM1[1723]<=16'd4790; ROM2[1723]<=16'd0; ROM3[1723]<=16'd23853; ROM4[1723]<=16'd57309;
ROM1[1724]<=16'd4816; ROM2[1724]<=16'd0; ROM3[1724]<=16'd23841; ROM4[1724]<=16'd57304;
ROM1[1725]<=16'd4836; ROM2[1725]<=16'd0; ROM3[1725]<=16'd23838; ROM4[1725]<=16'd57307;
ROM1[1726]<=16'd4829; ROM2[1726]<=16'd0; ROM3[1726]<=16'd23846; ROM4[1726]<=16'd57312;
ROM1[1727]<=16'd4803; ROM2[1727]<=16'd0; ROM3[1727]<=16'd23846; ROM4[1727]<=16'd57303;
ROM1[1728]<=16'd4789; ROM2[1728]<=16'd0; ROM3[1728]<=16'd23855; ROM4[1728]<=16'd57308;
ROM1[1729]<=16'd4777; ROM2[1729]<=16'd0; ROM3[1729]<=16'd23859; ROM4[1729]<=16'd57306;
ROM1[1730]<=16'd4761; ROM2[1730]<=16'd0; ROM3[1730]<=16'd23846; ROM4[1730]<=16'd57292;
ROM1[1731]<=16'd4772; ROM2[1731]<=16'd0; ROM3[1731]<=16'd23847; ROM4[1731]<=16'd57298;
ROM1[1732]<=16'd4799; ROM2[1732]<=16'd0; ROM3[1732]<=16'd23836; ROM4[1732]<=16'd57297;
ROM1[1733]<=16'd4831; ROM2[1733]<=16'd0; ROM3[1733]<=16'd23827; ROM4[1733]<=16'd57305;
ROM1[1734]<=16'd4831; ROM2[1734]<=16'd0; ROM3[1734]<=16'd23828; ROM4[1734]<=16'd57305;
ROM1[1735]<=16'd4809; ROM2[1735]<=16'd0; ROM3[1735]<=16'd23826; ROM4[1735]<=16'd57296;
ROM1[1736]<=16'd4793; ROM2[1736]<=16'd0; ROM3[1736]<=16'd23836; ROM4[1736]<=16'd57296;
ROM1[1737]<=16'd4789; ROM2[1737]<=16'd0; ROM3[1737]<=16'd23846; ROM4[1737]<=16'd57302;
ROM1[1738]<=16'd4779; ROM2[1738]<=16'd0; ROM3[1738]<=16'd23851; ROM4[1738]<=16'd57306;
ROM1[1739]<=16'd4772; ROM2[1739]<=16'd0; ROM3[1739]<=16'd23841; ROM4[1739]<=16'd57295;
ROM1[1740]<=16'd4798; ROM2[1740]<=16'd0; ROM3[1740]<=16'd23832; ROM4[1740]<=16'd57295;
ROM1[1741]<=16'd4825; ROM2[1741]<=16'd0; ROM3[1741]<=16'd23817; ROM4[1741]<=16'd57292;
ROM1[1742]<=16'd4821; ROM2[1742]<=16'd0; ROM3[1742]<=16'd23803; ROM4[1742]<=16'd57279;
ROM1[1743]<=16'd4805; ROM2[1743]<=16'd0; ROM3[1743]<=16'd23809; ROM4[1743]<=16'd57281;
ROM1[1744]<=16'd4784; ROM2[1744]<=16'd0; ROM3[1744]<=16'd23818; ROM4[1744]<=16'd57282;
ROM1[1745]<=16'd4777; ROM2[1745]<=16'd0; ROM3[1745]<=16'd23831; ROM4[1745]<=16'd57288;
ROM1[1746]<=16'd4787; ROM2[1746]<=16'd0; ROM3[1746]<=16'd23866; ROM4[1746]<=16'd57322;
ROM1[1747]<=16'd4810; ROM2[1747]<=16'd0; ROM3[1747]<=16'd23889; ROM4[1747]<=16'd57342;
ROM1[1748]<=16'd4802; ROM2[1748]<=16'd0; ROM3[1748]<=16'd23853; ROM4[1748]<=16'd57312;
ROM1[1749]<=16'd4787; ROM2[1749]<=16'd0; ROM3[1749]<=16'd23797; ROM4[1749]<=16'd57270;
ROM1[1750]<=16'd4782; ROM2[1750]<=16'd0; ROM3[1750]<=16'd23776; ROM4[1750]<=16'd57253;
ROM1[1751]<=16'd4767; ROM2[1751]<=16'd0; ROM3[1751]<=16'd23778; ROM4[1751]<=16'd57249;
ROM1[1752]<=16'd4763; ROM2[1752]<=16'd0; ROM3[1752]<=16'd23805; ROM4[1752]<=16'd57264;
ROM1[1753]<=16'd4757; ROM2[1753]<=16'd0; ROM3[1753]<=16'd23826; ROM4[1753]<=16'd57276;
ROM1[1754]<=16'd4733; ROM2[1754]<=16'd0; ROM3[1754]<=16'd23823; ROM4[1754]<=16'd57265;
ROM1[1755]<=16'd4709; ROM2[1755]<=16'd0; ROM3[1755]<=16'd23812; ROM4[1755]<=16'd57252;
ROM1[1756]<=16'd4713; ROM2[1756]<=16'd0; ROM3[1756]<=16'd23808; ROM4[1756]<=16'd57253;
ROM1[1757]<=16'd4748; ROM2[1757]<=16'd0; ROM3[1757]<=16'd23810; ROM4[1757]<=16'd57261;
ROM1[1758]<=16'd4770; ROM2[1758]<=16'd0; ROM3[1758]<=16'd23796; ROM4[1758]<=16'd57256;
ROM1[1759]<=16'd4765; ROM2[1759]<=16'd0; ROM3[1759]<=16'd23786; ROM4[1759]<=16'd57252;
ROM1[1760]<=16'd4773; ROM2[1760]<=16'd0; ROM3[1760]<=16'd23812; ROM4[1760]<=16'd57270;
ROM1[1761]<=16'd4769; ROM2[1761]<=16'd0; ROM3[1761]<=16'd23829; ROM4[1761]<=16'd57278;
ROM1[1762]<=16'd4754; ROM2[1762]<=16'd0; ROM3[1762]<=16'd23828; ROM4[1762]<=16'd57274;
ROM1[1763]<=16'd4746; ROM2[1763]<=16'd0; ROM3[1763]<=16'd23836; ROM4[1763]<=16'd57277;
ROM1[1764]<=16'd4750; ROM2[1764]<=16'd0; ROM3[1764]<=16'd23833; ROM4[1764]<=16'd57279;
ROM1[1765]<=16'd4775; ROM2[1765]<=16'd0; ROM3[1765]<=16'd23820; ROM4[1765]<=16'd57278;
ROM1[1766]<=16'd4808; ROM2[1766]<=16'd0; ROM3[1766]<=16'd23810; ROM4[1766]<=16'd57279;
ROM1[1767]<=16'd4809; ROM2[1767]<=16'd0; ROM3[1767]<=16'd23806; ROM4[1767]<=16'd57274;
ROM1[1768]<=16'd4776; ROM2[1768]<=16'd0; ROM3[1768]<=16'd23795; ROM4[1768]<=16'd57257;
ROM1[1769]<=16'd4757; ROM2[1769]<=16'd0; ROM3[1769]<=16'd23800; ROM4[1769]<=16'd57255;
ROM1[1770]<=16'd4754; ROM2[1770]<=16'd0; ROM3[1770]<=16'd23815; ROM4[1770]<=16'd57264;
ROM1[1771]<=16'd4754; ROM2[1771]<=16'd0; ROM3[1771]<=16'd23830; ROM4[1771]<=16'd57278;
ROM1[1772]<=16'd4761; ROM2[1772]<=16'd0; ROM3[1772]<=16'd23833; ROM4[1772]<=16'd57287;
ROM1[1773]<=16'd4784; ROM2[1773]<=16'd0; ROM3[1773]<=16'd23835; ROM4[1773]<=16'd57293;
ROM1[1774]<=16'd4817; ROM2[1774]<=16'd0; ROM3[1774]<=16'd23826; ROM4[1774]<=16'd57294;
ROM1[1775]<=16'd4830; ROM2[1775]<=16'd0; ROM3[1775]<=16'd23815; ROM4[1775]<=16'd57292;
ROM1[1776]<=16'd4825; ROM2[1776]<=16'd0; ROM3[1776]<=16'd23823; ROM4[1776]<=16'd57296;
ROM1[1777]<=16'd4807; ROM2[1777]<=16'd0; ROM3[1777]<=16'd23827; ROM4[1777]<=16'd57300;
ROM1[1778]<=16'd4795; ROM2[1778]<=16'd0; ROM3[1778]<=16'd23835; ROM4[1778]<=16'd57306;
ROM1[1779]<=16'd4781; ROM2[1779]<=16'd0; ROM3[1779]<=16'd23848; ROM4[1779]<=16'd57310;
ROM1[1780]<=16'd4765; ROM2[1780]<=16'd0; ROM3[1780]<=16'd23845; ROM4[1780]<=16'd57302;
ROM1[1781]<=16'd4779; ROM2[1781]<=16'd0; ROM3[1781]<=16'd23846; ROM4[1781]<=16'd57305;
ROM1[1782]<=16'd4818; ROM2[1782]<=16'd0; ROM3[1782]<=16'd23844; ROM4[1782]<=16'd57313;
ROM1[1783]<=16'd4836; ROM2[1783]<=16'd0; ROM3[1783]<=16'd23821; ROM4[1783]<=16'd57302;
ROM1[1784]<=16'd4825; ROM2[1784]<=16'd0; ROM3[1784]<=16'd23814; ROM4[1784]<=16'd57294;
ROM1[1785]<=16'd4809; ROM2[1785]<=16'd0; ROM3[1785]<=16'd23827; ROM4[1785]<=16'd57302;
ROM1[1786]<=16'd4794; ROM2[1786]<=16'd0; ROM3[1786]<=16'd23840; ROM4[1786]<=16'd57306;
ROM1[1787]<=16'd4793; ROM2[1787]<=16'd0; ROM3[1787]<=16'd23860; ROM4[1787]<=16'd57316;
ROM1[1788]<=16'd4778; ROM2[1788]<=16'd0; ROM3[1788]<=16'd23859; ROM4[1788]<=16'd57311;
ROM1[1789]<=16'd4764; ROM2[1789]<=16'd0; ROM3[1789]<=16'd23843; ROM4[1789]<=16'd57291;
ROM1[1790]<=16'd4795; ROM2[1790]<=16'd0; ROM3[1790]<=16'd23843; ROM4[1790]<=16'd57296;
ROM1[1791]<=16'd4837; ROM2[1791]<=16'd0; ROM3[1791]<=16'd23835; ROM4[1791]<=16'd57308;
ROM1[1792]<=16'd4819; ROM2[1792]<=16'd0; ROM3[1792]<=16'd23810; ROM4[1792]<=16'd57287;
ROM1[1793]<=16'd4787; ROM2[1793]<=16'd0; ROM3[1793]<=16'd23797; ROM4[1793]<=16'd57267;
ROM1[1794]<=16'd4764; ROM2[1794]<=16'd0; ROM3[1794]<=16'd23799; ROM4[1794]<=16'd57260;
ROM1[1795]<=16'd4744; ROM2[1795]<=16'd0; ROM3[1795]<=16'd23798; ROM4[1795]<=16'd57252;
ROM1[1796]<=16'd4745; ROM2[1796]<=16'd0; ROM3[1796]<=16'd23815; ROM4[1796]<=16'd57269;
ROM1[1797]<=16'd4749; ROM2[1797]<=16'd0; ROM3[1797]<=16'd23812; ROM4[1797]<=16'd57274;
ROM1[1798]<=16'd4751; ROM2[1798]<=16'd0; ROM3[1798]<=16'd23787; ROM4[1798]<=16'd57260;
ROM1[1799]<=16'd4782; ROM2[1799]<=16'd0; ROM3[1799]<=16'd23777; ROM4[1799]<=16'd57261;
ROM1[1800]<=16'd4807; ROM2[1800]<=16'd0; ROM3[1800]<=16'd23777; ROM4[1800]<=16'd57264;
ROM1[1801]<=16'd4805; ROM2[1801]<=16'd0; ROM3[1801]<=16'd23785; ROM4[1801]<=16'd57268;
ROM1[1802]<=16'd4782; ROM2[1802]<=16'd0; ROM3[1802]<=16'd23788; ROM4[1802]<=16'd57266;
ROM1[1803]<=16'd4765; ROM2[1803]<=16'd0; ROM3[1803]<=16'd23794; ROM4[1803]<=16'd57265;
ROM1[1804]<=16'd4757; ROM2[1804]<=16'd0; ROM3[1804]<=16'd23808; ROM4[1804]<=16'd57276;
ROM1[1805]<=16'd4752; ROM2[1805]<=16'd0; ROM3[1805]<=16'd23817; ROM4[1805]<=16'd57285;
ROM1[1806]<=16'd4781; ROM2[1806]<=16'd0; ROM3[1806]<=16'd23829; ROM4[1806]<=16'd57301;
ROM1[1807]<=16'd4816; ROM2[1807]<=16'd0; ROM3[1807]<=16'd23823; ROM4[1807]<=16'd57305;
ROM1[1808]<=16'd4816; ROM2[1808]<=16'd0; ROM3[1808]<=16'd23786; ROM4[1808]<=16'd57279;
ROM1[1809]<=16'd4796; ROM2[1809]<=16'd0; ROM3[1809]<=16'd23776; ROM4[1809]<=16'd57265;
ROM1[1810]<=16'd4775; ROM2[1810]<=16'd0; ROM3[1810]<=16'd23781; ROM4[1810]<=16'd57262;
ROM1[1811]<=16'd4753; ROM2[1811]<=16'd0; ROM3[1811]<=16'd23779; ROM4[1811]<=16'd57253;
ROM1[1812]<=16'd4747; ROM2[1812]<=16'd0; ROM3[1812]<=16'd23794; ROM4[1812]<=16'd57261;
ROM1[1813]<=16'd4742; ROM2[1813]<=16'd0; ROM3[1813]<=16'd23807; ROM4[1813]<=16'd57267;
ROM1[1814]<=16'd4748; ROM2[1814]<=16'd0; ROM3[1814]<=16'd23806; ROM4[1814]<=16'd57269;
ROM1[1815]<=16'd4786; ROM2[1815]<=16'd0; ROM3[1815]<=16'd23813; ROM4[1815]<=16'd57286;
ROM1[1816]<=16'd4835; ROM2[1816]<=16'd0; ROM3[1816]<=16'd23813; ROM4[1816]<=16'd57301;
ROM1[1817]<=16'd4838; ROM2[1817]<=16'd0; ROM3[1817]<=16'd23808; ROM4[1817]<=16'd57300;
ROM1[1818]<=16'd4794; ROM2[1818]<=16'd0; ROM3[1818]<=16'd23797; ROM4[1818]<=16'd57280;
ROM1[1819]<=16'd4756; ROM2[1819]<=16'd0; ROM3[1819]<=16'd23795; ROM4[1819]<=16'd57265;
ROM1[1820]<=16'd4745; ROM2[1820]<=16'd0; ROM3[1820]<=16'd23805; ROM4[1820]<=16'd57269;
ROM1[1821]<=16'd4733; ROM2[1821]<=16'd0; ROM3[1821]<=16'd23814; ROM4[1821]<=16'd57271;
ROM1[1822]<=16'd4742; ROM2[1822]<=16'd0; ROM3[1822]<=16'd23825; ROM4[1822]<=16'd57280;
ROM1[1823]<=16'd4760; ROM2[1823]<=16'd0; ROM3[1823]<=16'd23820; ROM4[1823]<=16'd57283;
ROM1[1824]<=16'd4788; ROM2[1824]<=16'd0; ROM3[1824]<=16'd23805; ROM4[1824]<=16'd57280;
ROM1[1825]<=16'd4812; ROM2[1825]<=16'd0; ROM3[1825]<=16'd23802; ROM4[1825]<=16'd57289;
ROM1[1826]<=16'd4803; ROM2[1826]<=16'd0; ROM3[1826]<=16'd23806; ROM4[1826]<=16'd57291;
ROM1[1827]<=16'd4780; ROM2[1827]<=16'd0; ROM3[1827]<=16'd23812; ROM4[1827]<=16'd57285;
ROM1[1828]<=16'd4772; ROM2[1828]<=16'd0; ROM3[1828]<=16'd23827; ROM4[1828]<=16'd57291;
ROM1[1829]<=16'd4765; ROM2[1829]<=16'd0; ROM3[1829]<=16'd23840; ROM4[1829]<=16'd57297;
ROM1[1830]<=16'd4745; ROM2[1830]<=16'd0; ROM3[1830]<=16'd23836; ROM4[1830]<=16'd57287;
ROM1[1831]<=16'd4750; ROM2[1831]<=16'd0; ROM3[1831]<=16'd23827; ROM4[1831]<=16'd57283;
ROM1[1832]<=16'd4776; ROM2[1832]<=16'd0; ROM3[1832]<=16'd23817; ROM4[1832]<=16'd57279;
ROM1[1833]<=16'd4791; ROM2[1833]<=16'd0; ROM3[1833]<=16'd23802; ROM4[1833]<=16'd57272;
ROM1[1834]<=16'd4795; ROM2[1834]<=16'd0; ROM3[1834]<=16'd23802; ROM4[1834]<=16'd57278;
ROM1[1835]<=16'd4787; ROM2[1835]<=16'd0; ROM3[1835]<=16'd23811; ROM4[1835]<=16'd57283;
ROM1[1836]<=16'd4772; ROM2[1836]<=16'd0; ROM3[1836]<=16'd23824; ROM4[1836]<=16'd57285;
ROM1[1837]<=16'd4757; ROM2[1837]<=16'd0; ROM3[1837]<=16'd23832; ROM4[1837]<=16'd57290;
ROM1[1838]<=16'd4743; ROM2[1838]<=16'd0; ROM3[1838]<=16'd23838; ROM4[1838]<=16'd57294;
ROM1[1839]<=16'd4741; ROM2[1839]<=16'd0; ROM3[1839]<=16'd23831; ROM4[1839]<=16'd57291;
ROM1[1840]<=16'd4769; ROM2[1840]<=16'd0; ROM3[1840]<=16'd23823; ROM4[1840]<=16'd57293;
ROM1[1841]<=16'd4808; ROM2[1841]<=16'd0; ROM3[1841]<=16'd23814; ROM4[1841]<=16'd57298;
ROM1[1842]<=16'd4815; ROM2[1842]<=16'd0; ROM3[1842]<=16'd23814; ROM4[1842]<=16'd57297;
ROM1[1843]<=16'd4791; ROM2[1843]<=16'd0; ROM3[1843]<=16'd23815; ROM4[1843]<=16'd57292;
ROM1[1844]<=16'd4767; ROM2[1844]<=16'd0; ROM3[1844]<=16'd23814; ROM4[1844]<=16'd57287;
ROM1[1845]<=16'd4751; ROM2[1845]<=16'd0; ROM3[1845]<=16'd23820; ROM4[1845]<=16'd57284;
ROM1[1846]<=16'd4731; ROM2[1846]<=16'd0; ROM3[1846]<=16'd23827; ROM4[1846]<=16'd57285;
ROM1[1847]<=16'd4735; ROM2[1847]<=16'd0; ROM3[1847]<=16'd23834; ROM4[1847]<=16'd57289;
ROM1[1848]<=16'd4747; ROM2[1848]<=16'd0; ROM3[1848]<=16'd23820; ROM4[1848]<=16'd57282;
ROM1[1849]<=16'd4773; ROM2[1849]<=16'd0; ROM3[1849]<=16'd23804; ROM4[1849]<=16'd57279;
ROM1[1850]<=16'd4797; ROM2[1850]<=16'd0; ROM3[1850]<=16'd23800; ROM4[1850]<=16'd57282;
ROM1[1851]<=16'd4781; ROM2[1851]<=16'd0; ROM3[1851]<=16'd23800; ROM4[1851]<=16'd57279;
ROM1[1852]<=16'd4755; ROM2[1852]<=16'd0; ROM3[1852]<=16'd23810; ROM4[1852]<=16'd57281;
ROM1[1853]<=16'd4754; ROM2[1853]<=16'd0; ROM3[1853]<=16'd23827; ROM4[1853]<=16'd57290;
ROM1[1854]<=16'd4749; ROM2[1854]<=16'd0; ROM3[1854]<=16'd23839; ROM4[1854]<=16'd57300;
ROM1[1855]<=16'd4742; ROM2[1855]<=16'd0; ROM3[1855]<=16'd23844; ROM4[1855]<=16'd57300;
ROM1[1856]<=16'd4762; ROM2[1856]<=16'd0; ROM3[1856]<=16'd23850; ROM4[1856]<=16'd57303;
ROM1[1857]<=16'd4792; ROM2[1857]<=16'd0; ROM3[1857]<=16'd23843; ROM4[1857]<=16'd57301;
ROM1[1858]<=16'd4813; ROM2[1858]<=16'd0; ROM3[1858]<=16'd23837; ROM4[1858]<=16'd57298;
ROM1[1859]<=16'd4817; ROM2[1859]<=16'd0; ROM3[1859]<=16'd23841; ROM4[1859]<=16'd57303;
ROM1[1860]<=16'd4796; ROM2[1860]<=16'd0; ROM3[1860]<=16'd23845; ROM4[1860]<=16'd57302;
ROM1[1861]<=16'd4776; ROM2[1861]<=16'd0; ROM3[1861]<=16'd23852; ROM4[1861]<=16'd57303;
ROM1[1862]<=16'd4750; ROM2[1862]<=16'd0; ROM3[1862]<=16'd23840; ROM4[1862]<=16'd57289;
ROM1[1863]<=16'd4720; ROM2[1863]<=16'd0; ROM3[1863]<=16'd23829; ROM4[1863]<=16'd57270;
ROM1[1864]<=16'd4725; ROM2[1864]<=16'd0; ROM3[1864]<=16'd23827; ROM4[1864]<=16'd57267;
ROM1[1865]<=16'd4754; ROM2[1865]<=16'd0; ROM3[1865]<=16'd23820; ROM4[1865]<=16'd57272;
ROM1[1866]<=16'd4791; ROM2[1866]<=16'd0; ROM3[1866]<=16'd23812; ROM4[1866]<=16'd57275;
ROM1[1867]<=16'd4789; ROM2[1867]<=16'd0; ROM3[1867]<=16'd23799; ROM4[1867]<=16'd57264;
ROM1[1868]<=16'd4774; ROM2[1868]<=16'd0; ROM3[1868]<=16'd23806; ROM4[1868]<=16'd57269;
ROM1[1869]<=16'd4768; ROM2[1869]<=16'd0; ROM3[1869]<=16'd23829; ROM4[1869]<=16'd57286;
ROM1[1870]<=16'd4742; ROM2[1870]<=16'd0; ROM3[1870]<=16'd23827; ROM4[1870]<=16'd57278;
ROM1[1871]<=16'd4737; ROM2[1871]<=16'd0; ROM3[1871]<=16'd23845; ROM4[1871]<=16'd57287;
ROM1[1872]<=16'd4746; ROM2[1872]<=16'd0; ROM3[1872]<=16'd23857; ROM4[1872]<=16'd57297;
ROM1[1873]<=16'd4721; ROM2[1873]<=16'd0; ROM3[1873]<=16'd23812; ROM4[1873]<=16'd57257;
ROM1[1874]<=16'd4745; ROM2[1874]<=16'd0; ROM3[1874]<=16'd23794; ROM4[1874]<=16'd57248;
ROM1[1875]<=16'd4766; ROM2[1875]<=16'd0; ROM3[1875]<=16'd23788; ROM4[1875]<=16'd57255;
ROM1[1876]<=16'd4743; ROM2[1876]<=16'd0; ROM3[1876]<=16'd23780; ROM4[1876]<=16'd57244;
ROM1[1877]<=16'd4728; ROM2[1877]<=16'd0; ROM3[1877]<=16'd23792; ROM4[1877]<=16'd57247;
ROM1[1878]<=16'd4722; ROM2[1878]<=16'd0; ROM3[1878]<=16'd23807; ROM4[1878]<=16'd57256;
ROM1[1879]<=16'd4710; ROM2[1879]<=16'd0; ROM3[1879]<=16'd23821; ROM4[1879]<=16'd57260;
ROM1[1880]<=16'd4703; ROM2[1880]<=16'd0; ROM3[1880]<=16'd23822; ROM4[1880]<=16'd57259;
ROM1[1881]<=16'd4718; ROM2[1881]<=16'd0; ROM3[1881]<=16'd23818; ROM4[1881]<=16'd57258;
ROM1[1882]<=16'd4746; ROM2[1882]<=16'd0; ROM3[1882]<=16'd23810; ROM4[1882]<=16'd57258;
ROM1[1883]<=16'd4772; ROM2[1883]<=16'd0; ROM3[1883]<=16'd23799; ROM4[1883]<=16'd57260;
ROM1[1884]<=16'd4762; ROM2[1884]<=16'd0; ROM3[1884]<=16'd23797; ROM4[1884]<=16'd57259;
ROM1[1885]<=16'd4744; ROM2[1885]<=16'd0; ROM3[1885]<=16'd23809; ROM4[1885]<=16'd57261;
ROM1[1886]<=16'd4726; ROM2[1886]<=16'd0; ROM3[1886]<=16'd23814; ROM4[1886]<=16'd57257;
ROM1[1887]<=16'd4712; ROM2[1887]<=16'd0; ROM3[1887]<=16'd23818; ROM4[1887]<=16'd57257;
ROM1[1888]<=16'd4709; ROM2[1888]<=16'd0; ROM3[1888]<=16'd23830; ROM4[1888]<=16'd57266;
ROM1[1889]<=16'd4718; ROM2[1889]<=16'd0; ROM3[1889]<=16'd23828; ROM4[1889]<=16'd57269;
ROM1[1890]<=16'd4746; ROM2[1890]<=16'd0; ROM3[1890]<=16'd23818; ROM4[1890]<=16'd57268;
ROM1[1891]<=16'd4787; ROM2[1891]<=16'd0; ROM3[1891]<=16'd23817; ROM4[1891]<=16'd57281;
ROM1[1892]<=16'd4793; ROM2[1892]<=16'd0; ROM3[1892]<=16'd23813; ROM4[1892]<=16'd57281;
ROM1[1893]<=16'd4778; ROM2[1893]<=16'd0; ROM3[1893]<=16'd23816; ROM4[1893]<=16'd57282;
ROM1[1894]<=16'd4772; ROM2[1894]<=16'd0; ROM3[1894]<=16'd23835; ROM4[1894]<=16'd57298;
ROM1[1895]<=16'd4765; ROM2[1895]<=16'd0; ROM3[1895]<=16'd23845; ROM4[1895]<=16'd57300;
ROM1[1896]<=16'd4749; ROM2[1896]<=16'd0; ROM3[1896]<=16'd23851; ROM4[1896]<=16'd57296;
ROM1[1897]<=16'd4760; ROM2[1897]<=16'd0; ROM3[1897]<=16'd23861; ROM4[1897]<=16'd57305;
ROM1[1898]<=16'd4774; ROM2[1898]<=16'd0; ROM3[1898]<=16'd23856; ROM4[1898]<=16'd57304;
ROM1[1899]<=16'd4793; ROM2[1899]<=16'd0; ROM3[1899]<=16'd23833; ROM4[1899]<=16'd57292;
ROM1[1900]<=16'd4815; ROM2[1900]<=16'd0; ROM3[1900]<=16'd23828; ROM4[1900]<=16'd57298;
ROM1[1901]<=16'd4799; ROM2[1901]<=16'd0; ROM3[1901]<=16'd23820; ROM4[1901]<=16'd57292;
ROM1[1902]<=16'd4773; ROM2[1902]<=16'd0; ROM3[1902]<=16'd23821; ROM4[1902]<=16'd57283;
ROM1[1903]<=16'd4763; ROM2[1903]<=16'd0; ROM3[1903]<=16'd23829; ROM4[1903]<=16'd57286;
ROM1[1904]<=16'd4748; ROM2[1904]<=16'd0; ROM3[1904]<=16'd23835; ROM4[1904]<=16'd57287;
ROM1[1905]<=16'd4740; ROM2[1905]<=16'd0; ROM3[1905]<=16'd23843; ROM4[1905]<=16'd57288;
ROM1[1906]<=16'd4753; ROM2[1906]<=16'd0; ROM3[1906]<=16'd23839; ROM4[1906]<=16'd57287;
ROM1[1907]<=16'd4780; ROM2[1907]<=16'd0; ROM3[1907]<=16'd23825; ROM4[1907]<=16'd57284;
ROM1[1908]<=16'd4807; ROM2[1908]<=16'd0; ROM3[1908]<=16'd23816; ROM4[1908]<=16'd57284;
ROM1[1909]<=16'd4803; ROM2[1909]<=16'd0; ROM3[1909]<=16'd23818; ROM4[1909]<=16'd57286;
ROM1[1910]<=16'd4793; ROM2[1910]<=16'd0; ROM3[1910]<=16'd23831; ROM4[1910]<=16'd57298;
ROM1[1911]<=16'd4787; ROM2[1911]<=16'd0; ROM3[1911]<=16'd23847; ROM4[1911]<=16'd57308;
ROM1[1912]<=16'd4756; ROM2[1912]<=16'd0; ROM3[1912]<=16'd23842; ROM4[1912]<=16'd57294;
ROM1[1913]<=16'd4740; ROM2[1913]<=16'd0; ROM3[1913]<=16'd23843; ROM4[1913]<=16'd57288;
ROM1[1914]<=16'd4752; ROM2[1914]<=16'd0; ROM3[1914]<=16'd23847; ROM4[1914]<=16'd57294;
ROM1[1915]<=16'd4785; ROM2[1915]<=16'd0; ROM3[1915]<=16'd23845; ROM4[1915]<=16'd57301;
ROM1[1916]<=16'd4809; ROM2[1916]<=16'd0; ROM3[1916]<=16'd23826; ROM4[1916]<=16'd57290;
ROM1[1917]<=16'd4791; ROM2[1917]<=16'd0; ROM3[1917]<=16'd23803; ROM4[1917]<=16'd57271;
ROM1[1918]<=16'd4783; ROM2[1918]<=16'd0; ROM3[1918]<=16'd23818; ROM4[1918]<=16'd57281;
ROM1[1919]<=16'd4769; ROM2[1919]<=16'd0; ROM3[1919]<=16'd23836; ROM4[1919]<=16'd57289;
ROM1[1920]<=16'd4747; ROM2[1920]<=16'd0; ROM3[1920]<=16'd23833; ROM4[1920]<=16'd57284;
ROM1[1921]<=16'd4741; ROM2[1921]<=16'd0; ROM3[1921]<=16'd23846; ROM4[1921]<=16'd57291;
ROM1[1922]<=16'd4744; ROM2[1922]<=16'd0; ROM3[1922]<=16'd23852; ROM4[1922]<=16'd57296;
ROM1[1923]<=16'd4752; ROM2[1923]<=16'd0; ROM3[1923]<=16'd23839; ROM4[1923]<=16'd57287;
ROM1[1924]<=16'd4782; ROM2[1924]<=16'd0; ROM3[1924]<=16'd23826; ROM4[1924]<=16'd57286;
ROM1[1925]<=16'd4808; ROM2[1925]<=16'd0; ROM3[1925]<=16'd23825; ROM4[1925]<=16'd57295;
ROM1[1926]<=16'd4780; ROM2[1926]<=16'd0; ROM3[1926]<=16'd23811; ROM4[1926]<=16'd57278;
ROM1[1927]<=16'd4744; ROM2[1927]<=16'd0; ROM3[1927]<=16'd23796; ROM4[1927]<=16'd57262;
ROM1[1928]<=16'd4740; ROM2[1928]<=16'd0; ROM3[1928]<=16'd23816; ROM4[1928]<=16'd57275;
ROM1[1929]<=16'd4721; ROM2[1929]<=16'd0; ROM3[1929]<=16'd23825; ROM4[1929]<=16'd57277;
ROM1[1930]<=16'd4706; ROM2[1930]<=16'd0; ROM3[1930]<=16'd23813; ROM4[1930]<=16'd57268;
ROM1[1931]<=16'd4716; ROM2[1931]<=16'd0; ROM3[1931]<=16'd23804; ROM4[1931]<=16'd57261;
ROM1[1932]<=16'd4754; ROM2[1932]<=16'd0; ROM3[1932]<=16'd23797; ROM4[1932]<=16'd57262;
ROM1[1933]<=16'd4789; ROM2[1933]<=16'd0; ROM3[1933]<=16'd23792; ROM4[1933]<=16'd57267;
ROM1[1934]<=16'd4789; ROM2[1934]<=16'd0; ROM3[1934]<=16'd23797; ROM4[1934]<=16'd57272;
ROM1[1935]<=16'd4778; ROM2[1935]<=16'd0; ROM3[1935]<=16'd23813; ROM4[1935]<=16'd57279;
ROM1[1936]<=16'd4769; ROM2[1936]<=16'd0; ROM3[1936]<=16'd23834; ROM4[1936]<=16'd57290;
ROM1[1937]<=16'd4769; ROM2[1937]<=16'd0; ROM3[1937]<=16'd23851; ROM4[1937]<=16'd57302;
ROM1[1938]<=16'd4771; ROM2[1938]<=16'd0; ROM3[1938]<=16'd23871; ROM4[1938]<=16'd57318;
ROM1[1939]<=16'd4770; ROM2[1939]<=16'd0; ROM3[1939]<=16'd23866; ROM4[1939]<=16'd57311;
ROM1[1940]<=16'd4787; ROM2[1940]<=16'd0; ROM3[1940]<=16'd23843; ROM4[1940]<=16'd57301;
ROM1[1941]<=16'd4811; ROM2[1941]<=16'd0; ROM3[1941]<=16'd23823; ROM4[1941]<=16'd57298;
ROM1[1942]<=16'd4803; ROM2[1942]<=16'd0; ROM3[1942]<=16'd23814; ROM4[1942]<=16'd57290;
ROM1[1943]<=16'd4790; ROM2[1943]<=16'd0; ROM3[1943]<=16'd23828; ROM4[1943]<=16'd57295;
ROM1[1944]<=16'd4784; ROM2[1944]<=16'd0; ROM3[1944]<=16'd23844; ROM4[1944]<=16'd57302;
ROM1[1945]<=16'd4778; ROM2[1945]<=16'd0; ROM3[1945]<=16'd23857; ROM4[1945]<=16'd57309;
ROM1[1946]<=16'd4769; ROM2[1946]<=16'd0; ROM3[1946]<=16'd23871; ROM4[1946]<=16'd57315;
ROM1[1947]<=16'd4764; ROM2[1947]<=16'd0; ROM3[1947]<=16'd23871; ROM4[1947]<=16'd57316;
ROM1[1948]<=16'd4774; ROM2[1948]<=16'd0; ROM3[1948]<=16'd23856; ROM4[1948]<=16'd57310;
ROM1[1949]<=16'd4797; ROM2[1949]<=16'd0; ROM3[1949]<=16'd23833; ROM4[1949]<=16'd57303;
ROM1[1950]<=16'd4817; ROM2[1950]<=16'd0; ROM3[1950]<=16'd23822; ROM4[1950]<=16'd57298;
ROM1[1951]<=16'd4812; ROM2[1951]<=16'd0; ROM3[1951]<=16'd23825; ROM4[1951]<=16'd57298;
ROM1[1952]<=16'd4796; ROM2[1952]<=16'd0; ROM3[1952]<=16'd23840; ROM4[1952]<=16'd57306;
ROM1[1953]<=16'd4796; ROM2[1953]<=16'd0; ROM3[1953]<=16'd23861; ROM4[1953]<=16'd57315;
ROM1[1954]<=16'd4789; ROM2[1954]<=16'd0; ROM3[1954]<=16'd23875; ROM4[1954]<=16'd57322;
ROM1[1955]<=16'd4773; ROM2[1955]<=16'd0; ROM3[1955]<=16'd23867; ROM4[1955]<=16'd57316;
ROM1[1956]<=16'd4762; ROM2[1956]<=16'd0; ROM3[1956]<=16'd23840; ROM4[1956]<=16'd57292;
ROM1[1957]<=16'd4778; ROM2[1957]<=16'd0; ROM3[1957]<=16'd23818; ROM4[1957]<=16'd57283;
ROM1[1958]<=16'd4790; ROM2[1958]<=16'd0; ROM3[1958]<=16'd23792; ROM4[1958]<=16'd57269;
ROM1[1959]<=16'd4795; ROM2[1959]<=16'd0; ROM3[1959]<=16'd23796; ROM4[1959]<=16'd57274;
ROM1[1960]<=16'd4801; ROM2[1960]<=16'd0; ROM3[1960]<=16'd23824; ROM4[1960]<=16'd57300;
ROM1[1961]<=16'd4783; ROM2[1961]<=16'd0; ROM3[1961]<=16'd23828; ROM4[1961]<=16'd57296;
ROM1[1962]<=16'd4756; ROM2[1962]<=16'd0; ROM3[1962]<=16'd23821; ROM4[1962]<=16'd57288;
ROM1[1963]<=16'd4744; ROM2[1963]<=16'd0; ROM3[1963]<=16'd23829; ROM4[1963]<=16'd57288;
ROM1[1964]<=16'd4754; ROM2[1964]<=16'd0; ROM3[1964]<=16'd23831; ROM4[1964]<=16'd57289;
ROM1[1965]<=16'd4785; ROM2[1965]<=16'd0; ROM3[1965]<=16'd23826; ROM4[1965]<=16'd57295;
ROM1[1966]<=16'd4814; ROM2[1966]<=16'd0; ROM3[1966]<=16'd23809; ROM4[1966]<=16'd57291;
ROM1[1967]<=16'd4803; ROM2[1967]<=16'd0; ROM3[1967]<=16'd23789; ROM4[1967]<=16'd57275;
ROM1[1968]<=16'd4777; ROM2[1968]<=16'd0; ROM3[1968]<=16'd23788; ROM4[1968]<=16'd57265;
ROM1[1969]<=16'd4757; ROM2[1969]<=16'd0; ROM3[1969]<=16'd23793; ROM4[1969]<=16'd57262;
ROM1[1970]<=16'd4756; ROM2[1970]<=16'd0; ROM3[1970]<=16'd23806; ROM4[1970]<=16'd57273;
ROM1[1971]<=16'd4747; ROM2[1971]<=16'd0; ROM3[1971]<=16'd23817; ROM4[1971]<=16'd57279;
ROM1[1972]<=16'd4730; ROM2[1972]<=16'd0; ROM3[1972]<=16'd23802; ROM4[1972]<=16'd57265;
ROM1[1973]<=16'd4737; ROM2[1973]<=16'd0; ROM3[1973]<=16'd23786; ROM4[1973]<=16'd57256;
ROM1[1974]<=16'd4769; ROM2[1974]<=16'd0; ROM3[1974]<=16'd23780; ROM4[1974]<=16'd57258;
ROM1[1975]<=16'd4788; ROM2[1975]<=16'd0; ROM3[1975]<=16'd23780; ROM4[1975]<=16'd57267;
ROM1[1976]<=16'd4777; ROM2[1976]<=16'd0; ROM3[1976]<=16'd23784; ROM4[1976]<=16'd57268;
ROM1[1977]<=16'd4750; ROM2[1977]<=16'd0; ROM3[1977]<=16'd23790; ROM4[1977]<=16'd57257;
ROM1[1978]<=16'd4745; ROM2[1978]<=16'd0; ROM3[1978]<=16'd23804; ROM4[1978]<=16'd57267;
ROM1[1979]<=16'd4739; ROM2[1979]<=16'd0; ROM3[1979]<=16'd23816; ROM4[1979]<=16'd57277;
ROM1[1980]<=16'd4719; ROM2[1980]<=16'd0; ROM3[1980]<=16'd23806; ROM4[1980]<=16'd57268;
ROM1[1981]<=16'd4735; ROM2[1981]<=16'd0; ROM3[1981]<=16'd23803; ROM4[1981]<=16'd57269;
ROM1[1982]<=16'd4779; ROM2[1982]<=16'd0; ROM3[1982]<=16'd23810; ROM4[1982]<=16'd57279;
ROM1[1983]<=16'd4819; ROM2[1983]<=16'd0; ROM3[1983]<=16'd23810; ROM4[1983]<=16'd57290;
ROM1[1984]<=16'd4814; ROM2[1984]<=16'd0; ROM3[1984]<=16'd23813; ROM4[1984]<=16'd57290;
ROM1[1985]<=16'd4781; ROM2[1985]<=16'd0; ROM3[1985]<=16'd23805; ROM4[1985]<=16'd57276;
ROM1[1986]<=16'd4755; ROM2[1986]<=16'd0; ROM3[1986]<=16'd23804; ROM4[1986]<=16'd57268;
ROM1[1987]<=16'd4721; ROM2[1987]<=16'd0; ROM3[1987]<=16'd23793; ROM4[1987]<=16'd57245;
ROM1[1988]<=16'd4719; ROM2[1988]<=16'd0; ROM3[1988]<=16'd23797; ROM4[1988]<=16'd57247;
ROM1[1989]<=16'd4735; ROM2[1989]<=16'd0; ROM3[1989]<=16'd23802; ROM4[1989]<=16'd57256;
ROM1[1990]<=16'd4748; ROM2[1990]<=16'd0; ROM3[1990]<=16'd23780; ROM4[1990]<=16'd57245;
ROM1[1991]<=16'd4777; ROM2[1991]<=16'd0; ROM3[1991]<=16'd23769; ROM4[1991]<=16'd57245;
ROM1[1992]<=16'd4783; ROM2[1992]<=16'd0; ROM3[1992]<=16'd23770; ROM4[1992]<=16'd57245;
ROM1[1993]<=16'd4772; ROM2[1993]<=16'd0; ROM3[1993]<=16'd23779; ROM4[1993]<=16'd57252;
ROM1[1994]<=16'd4756; ROM2[1994]<=16'd0; ROM3[1994]<=16'd23794; ROM4[1994]<=16'd57257;
ROM1[1995]<=16'd4750; ROM2[1995]<=16'd0; ROM3[1995]<=16'd23810; ROM4[1995]<=16'd57264;
ROM1[1996]<=16'd4762; ROM2[1996]<=16'd0; ROM3[1996]<=16'd23837; ROM4[1996]<=16'd57288;
ROM1[1997]<=16'd4757; ROM2[1997]<=16'd0; ROM3[1997]<=16'd23838; ROM4[1997]<=16'd57285;
ROM1[1998]<=16'd4752; ROM2[1998]<=16'd0; ROM3[1998]<=16'd23805; ROM4[1998]<=16'd57258;
ROM1[1999]<=16'd4786; ROM2[1999]<=16'd0; ROM3[1999]<=16'd23790; ROM4[1999]<=16'd57259;
ROM1[2000]<=16'd4807; ROM2[2000]<=16'd0; ROM3[2000]<=16'd23796; ROM4[2000]<=16'd57274;
ROM1[2001]<=16'd4802; ROM2[2001]<=16'd0; ROM3[2001]<=16'd23808; ROM4[2001]<=16'd57279;
ROM1[2002]<=16'd4779; ROM2[2002]<=16'd0; ROM3[2002]<=16'd23807; ROM4[2002]<=16'd57272;
ROM1[2003]<=16'd4756; ROM2[2003]<=16'd0; ROM3[2003]<=16'd23807; ROM4[2003]<=16'd57269;
ROM1[2004]<=16'd4726; ROM2[2004]<=16'd0; ROM3[2004]<=16'd23798; ROM4[2004]<=16'd57251;
ROM1[2005]<=16'd4712; ROM2[2005]<=16'd0; ROM3[2005]<=16'd23790; ROM4[2005]<=16'd57240;
ROM1[2006]<=16'd4736; ROM2[2006]<=16'd0; ROM3[2006]<=16'd23798; ROM4[2006]<=16'd57255;
ROM1[2007]<=16'd4774; ROM2[2007]<=16'd0; ROM3[2007]<=16'd23795; ROM4[2007]<=16'd57263;
ROM1[2008]<=16'd4801; ROM2[2008]<=16'd0; ROM3[2008]<=16'd23787; ROM4[2008]<=16'd57266;
ROM1[2009]<=16'd4792; ROM2[2009]<=16'd0; ROM3[2009]<=16'd23791; ROM4[2009]<=16'd57270;
ROM1[2010]<=16'd4768; ROM2[2010]<=16'd0; ROM3[2010]<=16'd23793; ROM4[2010]<=16'd57264;
ROM1[2011]<=16'd4741; ROM2[2011]<=16'd0; ROM3[2011]<=16'd23791; ROM4[2011]<=16'd57255;
ROM1[2012]<=16'd4720; ROM2[2012]<=16'd0; ROM3[2012]<=16'd23791; ROM4[2012]<=16'd57252;
ROM1[2013]<=16'd4712; ROM2[2013]<=16'd0; ROM3[2013]<=16'd23800; ROM4[2013]<=16'd57260;
ROM1[2014]<=16'd4722; ROM2[2014]<=16'd0; ROM3[2014]<=16'd23806; ROM4[2014]<=16'd57269;
ROM1[2015]<=16'd4749; ROM2[2015]<=16'd0; ROM3[2015]<=16'd23801; ROM4[2015]<=16'd57271;
ROM1[2016]<=16'd4783; ROM2[2016]<=16'd0; ROM3[2016]<=16'd23790; ROM4[2016]<=16'd57271;
ROM1[2017]<=16'd4790; ROM2[2017]<=16'd0; ROM3[2017]<=16'd23789; ROM4[2017]<=16'd57273;
ROM1[2018]<=16'd4778; ROM2[2018]<=16'd0; ROM3[2018]<=16'd23799; ROM4[2018]<=16'd57276;
ROM1[2019]<=16'd4762; ROM2[2019]<=16'd0; ROM3[2019]<=16'd23806; ROM4[2019]<=16'd57276;
ROM1[2020]<=16'd4745; ROM2[2020]<=16'd0; ROM3[2020]<=16'd23808; ROM4[2020]<=16'd57271;
ROM1[2021]<=16'd4729; ROM2[2021]<=16'd0; ROM3[2021]<=16'd23813; ROM4[2021]<=16'd57268;
ROM1[2022]<=16'd4733; ROM2[2022]<=16'd0; ROM3[2022]<=16'd23813; ROM4[2022]<=16'd57272;
ROM1[2023]<=16'd4753; ROM2[2023]<=16'd0; ROM3[2023]<=16'd23807; ROM4[2023]<=16'd57272;
ROM1[2024]<=16'd4788; ROM2[2024]<=16'd0; ROM3[2024]<=16'd23800; ROM4[2024]<=16'd57274;
ROM1[2025]<=16'd4801; ROM2[2025]<=16'd0; ROM3[2025]<=16'd23788; ROM4[2025]<=16'd57270;
ROM1[2026]<=16'd4782; ROM2[2026]<=16'd0; ROM3[2026]<=16'd23783; ROM4[2026]<=16'd57264;
ROM1[2027]<=16'd4770; ROM2[2027]<=16'd0; ROM3[2027]<=16'd23797; ROM4[2027]<=16'd57270;
ROM1[2028]<=16'd4773; ROM2[2028]<=16'd0; ROM3[2028]<=16'd23823; ROM4[2028]<=16'd57289;
ROM1[2029]<=16'd4775; ROM2[2029]<=16'd0; ROM3[2029]<=16'd23845; ROM4[2029]<=16'd57304;
ROM1[2030]<=16'd4756; ROM2[2030]<=16'd0; ROM3[2030]<=16'd23838; ROM4[2030]<=16'd57295;
ROM1[2031]<=16'd4756; ROM2[2031]<=16'd0; ROM3[2031]<=16'd23825; ROM4[2031]<=16'd57286;
ROM1[2032]<=16'd4787; ROM2[2032]<=16'd0; ROM3[2032]<=16'd23815; ROM4[2032]<=16'd57285;
ROM1[2033]<=16'd4808; ROM2[2033]<=16'd0; ROM3[2033]<=16'd23795; ROM4[2033]<=16'd57279;
ROM1[2034]<=16'd4807; ROM2[2034]<=16'd0; ROM3[2034]<=16'd23803; ROM4[2034]<=16'd57285;
ROM1[2035]<=16'd4799; ROM2[2035]<=16'd0; ROM3[2035]<=16'd23819; ROM4[2035]<=16'd57295;
ROM1[2036]<=16'd4785; ROM2[2036]<=16'd0; ROM3[2036]<=16'd23825; ROM4[2036]<=16'd57299;
ROM1[2037]<=16'd4773; ROM2[2037]<=16'd0; ROM3[2037]<=16'd23836; ROM4[2037]<=16'd57301;
ROM1[2038]<=16'd4756; ROM2[2038]<=16'd0; ROM3[2038]<=16'd23828; ROM4[2038]<=16'd57292;
ROM1[2039]<=16'd4744; ROM2[2039]<=16'd0; ROM3[2039]<=16'd23807; ROM4[2039]<=16'd57269;
ROM1[2040]<=16'd4754; ROM2[2040]<=16'd0; ROM3[2040]<=16'd23785; ROM4[2040]<=16'd57251;
ROM1[2041]<=16'd4789; ROM2[2041]<=16'd0; ROM3[2041]<=16'd23781; ROM4[2041]<=16'd57260;
ROM1[2042]<=16'd4827; ROM2[2042]<=16'd0; ROM3[2042]<=16'd23814; ROM4[2042]<=16'd57293;
ROM1[2043]<=16'd4815; ROM2[2043]<=16'd0; ROM3[2043]<=16'd23825; ROM4[2043]<=16'd57297;
ROM1[2044]<=16'd4763; ROM2[2044]<=16'd0; ROM3[2044]<=16'd23802; ROM4[2044]<=16'd57270;
ROM1[2045]<=16'd4734; ROM2[2045]<=16'd0; ROM3[2045]<=16'd23793; ROM4[2045]<=16'd57254;
ROM1[2046]<=16'd4710; ROM2[2046]<=16'd0; ROM3[2046]<=16'd23795; ROM4[2046]<=16'd57246;
ROM1[2047]<=16'd4711; ROM2[2047]<=16'd0; ROM3[2047]<=16'd23800; ROM4[2047]<=16'd57249;
ROM1[2048]<=16'd4747; ROM2[2048]<=16'd0; ROM3[2048]<=16'd23804; ROM4[2048]<=16'd57262;
ROM1[2049]<=16'd4789; ROM2[2049]<=16'd0; ROM3[2049]<=16'd23795; ROM4[2049]<=16'd57265;
ROM1[2050]<=16'd4793; ROM2[2050]<=16'd0; ROM3[2050]<=16'd23776; ROM4[2050]<=16'd57254;
ROM1[2051]<=16'd4780; ROM2[2051]<=16'd0; ROM3[2051]<=16'd23778; ROM4[2051]<=16'd57252;
ROM1[2052]<=16'd4767; ROM2[2052]<=16'd0; ROM3[2052]<=16'd23790; ROM4[2052]<=16'd57259;
ROM1[2053]<=16'd4754; ROM2[2053]<=16'd0; ROM3[2053]<=16'd23800; ROM4[2053]<=16'd57261;
ROM1[2054]<=16'd4740; ROM2[2054]<=16'd0; ROM3[2054]<=16'd23806; ROM4[2054]<=16'd57260;
ROM1[2055]<=16'd4736; ROM2[2055]<=16'd0; ROM3[2055]<=16'd23807; ROM4[2055]<=16'd57258;
ROM1[2056]<=16'd4755; ROM2[2056]<=16'd0; ROM3[2056]<=16'd23809; ROM4[2056]<=16'd57267;
ROM1[2057]<=16'd4783; ROM2[2057]<=16'd0; ROM3[2057]<=16'd23793; ROM4[2057]<=16'd57265;
ROM1[2058]<=16'd4802; ROM2[2058]<=16'd0; ROM3[2058]<=16'd23772; ROM4[2058]<=16'd57257;
ROM1[2059]<=16'd4798; ROM2[2059]<=16'd0; ROM3[2059]<=16'd23773; ROM4[2059]<=16'd57259;
ROM1[2060]<=16'd4784; ROM2[2060]<=16'd0; ROM3[2060]<=16'd23781; ROM4[2060]<=16'd57262;
ROM1[2061]<=16'd4776; ROM2[2061]<=16'd0; ROM3[2061]<=16'd23798; ROM4[2061]<=16'd57271;
ROM1[2062]<=16'd4774; ROM2[2062]<=16'd0; ROM3[2062]<=16'd23817; ROM4[2062]<=16'd57285;
ROM1[2063]<=16'd4749; ROM2[2063]<=16'd0; ROM3[2063]<=16'd23812; ROM4[2063]<=16'd57276;
ROM1[2064]<=16'd4745; ROM2[2064]<=16'd0; ROM3[2064]<=16'd23802; ROM4[2064]<=16'd57269;
ROM1[2065]<=16'd4766; ROM2[2065]<=16'd0; ROM3[2065]<=16'd23789; ROM4[2065]<=16'd57262;
ROM1[2066]<=16'd4801; ROM2[2066]<=16'd0; ROM3[2066]<=16'd23785; ROM4[2066]<=16'd57268;
ROM1[2067]<=16'd4811; ROM2[2067]<=16'd0; ROM3[2067]<=16'd23790; ROM4[2067]<=16'd57279;
ROM1[2068]<=16'd4788; ROM2[2068]<=16'd0; ROM3[2068]<=16'd23788; ROM4[2068]<=16'd57274;
ROM1[2069]<=16'd4770; ROM2[2069]<=16'd0; ROM3[2069]<=16'd23795; ROM4[2069]<=16'd57275;
ROM1[2070]<=16'd4758; ROM2[2070]<=16'd0; ROM3[2070]<=16'd23800; ROM4[2070]<=16'd57275;
ROM1[2071]<=16'd4751; ROM2[2071]<=16'd0; ROM3[2071]<=16'd23809; ROM4[2071]<=16'd57276;
ROM1[2072]<=16'd4751; ROM2[2072]<=16'd0; ROM3[2072]<=16'd23807; ROM4[2072]<=16'd57270;
ROM1[2073]<=16'd4767; ROM2[2073]<=16'd0; ROM3[2073]<=16'd23797; ROM4[2073]<=16'd57269;
ROM1[2074]<=16'd4792; ROM2[2074]<=16'd0; ROM3[2074]<=16'd23783; ROM4[2074]<=16'd57267;
ROM1[2075]<=16'd4803; ROM2[2075]<=16'd0; ROM3[2075]<=16'd23775; ROM4[2075]<=16'd57267;
ROM1[2076]<=16'd4795; ROM2[2076]<=16'd0; ROM3[2076]<=16'd23787; ROM4[2076]<=16'd57272;
ROM1[2077]<=16'd4767; ROM2[2077]<=16'd0; ROM3[2077]<=16'd23788; ROM4[2077]<=16'd57262;
ROM1[2078]<=16'd4748; ROM2[2078]<=16'd0; ROM3[2078]<=16'd23793; ROM4[2078]<=16'd57260;
ROM1[2079]<=16'd4733; ROM2[2079]<=16'd0; ROM3[2079]<=16'd23796; ROM4[2079]<=16'd57260;
ROM1[2080]<=16'd4729; ROM2[2080]<=16'd0; ROM3[2080]<=16'd23800; ROM4[2080]<=16'd57264;
ROM1[2081]<=16'd4744; ROM2[2081]<=16'd0; ROM3[2081]<=16'd23804; ROM4[2081]<=16'd57271;
ROM1[2082]<=16'd4771; ROM2[2082]<=16'd0; ROM3[2082]<=16'd23791; ROM4[2082]<=16'd57266;
ROM1[2083]<=16'd4792; ROM2[2083]<=16'd0; ROM3[2083]<=16'd23783; ROM4[2083]<=16'd57266;
ROM1[2084]<=16'd4787; ROM2[2084]<=16'd0; ROM3[2084]<=16'd23790; ROM4[2084]<=16'd57272;
ROM1[2085]<=16'd4771; ROM2[2085]<=16'd0; ROM3[2085]<=16'd23799; ROM4[2085]<=16'd57275;
ROM1[2086]<=16'd4773; ROM2[2086]<=16'd0; ROM3[2086]<=16'd23821; ROM4[2086]<=16'd57287;
ROM1[2087]<=16'd4789; ROM2[2087]<=16'd0; ROM3[2087]<=16'd23858; ROM4[2087]<=16'd57319;
ROM1[2088]<=16'd4788; ROM2[2088]<=16'd0; ROM3[2088]<=16'd23874; ROM4[2088]<=16'd57330;
ROM1[2089]<=16'd4769; ROM2[2089]<=16'd0; ROM3[2089]<=16'd23847; ROM4[2089]<=16'd57304;
ROM1[2090]<=16'd4760; ROM2[2090]<=16'd0; ROM3[2090]<=16'd23804; ROM4[2090]<=16'd57273;
ROM1[2091]<=16'd4766; ROM2[2091]<=16'd0; ROM3[2091]<=16'd23763; ROM4[2091]<=16'd57247;
ROM1[2092]<=16'd4754; ROM2[2092]<=16'd0; ROM3[2092]<=16'd23746; ROM4[2092]<=16'd57231;
ROM1[2093]<=16'd4755; ROM2[2093]<=16'd0; ROM3[2093]<=16'd23770; ROM4[2093]<=16'd57250;
ROM1[2094]<=16'd4751; ROM2[2094]<=16'd0; ROM3[2094]<=16'd23797; ROM4[2094]<=16'd57269;
ROM1[2095]<=16'd4734; ROM2[2095]<=16'd0; ROM3[2095]<=16'd23805; ROM4[2095]<=16'd57268;
ROM1[2096]<=16'd4716; ROM2[2096]<=16'd0; ROM3[2096]<=16'd23805; ROM4[2096]<=16'd57261;
ROM1[2097]<=16'd4717; ROM2[2097]<=16'd0; ROM3[2097]<=16'd23800; ROM4[2097]<=16'd57255;
ROM1[2098]<=16'd4742; ROM2[2098]<=16'd0; ROM3[2098]<=16'd23795; ROM4[2098]<=16'd57255;
ROM1[2099]<=16'd4783; ROM2[2099]<=16'd0; ROM3[2099]<=16'd23788; ROM4[2099]<=16'd57262;
ROM1[2100]<=16'd4806; ROM2[2100]<=16'd0; ROM3[2100]<=16'd23790; ROM4[2100]<=16'd57272;
ROM1[2101]<=16'd4792; ROM2[2101]<=16'd0; ROM3[2101]<=16'd23796; ROM4[2101]<=16'd57278;
ROM1[2102]<=16'd4767; ROM2[2102]<=16'd0; ROM3[2102]<=16'd23793; ROM4[2102]<=16'd57272;
ROM1[2103]<=16'd4758; ROM2[2103]<=16'd0; ROM3[2103]<=16'd23806; ROM4[2103]<=16'd57274;
ROM1[2104]<=16'd4763; ROM2[2104]<=16'd0; ROM3[2104]<=16'd23834; ROM4[2104]<=16'd57294;
ROM1[2105]<=16'd4752; ROM2[2105]<=16'd0; ROM3[2105]<=16'd23832; ROM4[2105]<=16'd57284;
ROM1[2106]<=16'd4755; ROM2[2106]<=16'd0; ROM3[2106]<=16'd23824; ROM4[2106]<=16'd57278;
ROM1[2107]<=16'd4786; ROM2[2107]<=16'd0; ROM3[2107]<=16'd23812; ROM4[2107]<=16'd57277;
ROM1[2108]<=16'd4795; ROM2[2108]<=16'd0; ROM3[2108]<=16'd23783; ROM4[2108]<=16'd57259;
ROM1[2109]<=16'd4792; ROM2[2109]<=16'd0; ROM3[2109]<=16'd23786; ROM4[2109]<=16'd57263;
ROM1[2110]<=16'd4785; ROM2[2110]<=16'd0; ROM3[2110]<=16'd23805; ROM4[2110]<=16'd57274;
ROM1[2111]<=16'd4760; ROM2[2111]<=16'd0; ROM3[2111]<=16'd23806; ROM4[2111]<=16'd57265;
ROM1[2112]<=16'd4753; ROM2[2112]<=16'd0; ROM3[2112]<=16'd23817; ROM4[2112]<=16'd57273;
ROM1[2113]<=16'd4759; ROM2[2113]<=16'd0; ROM3[2113]<=16'd23834; ROM4[2113]<=16'd57290;
ROM1[2114]<=16'd4755; ROM2[2114]<=16'd0; ROM3[2114]<=16'd23817; ROM4[2114]<=16'd57278;
ROM1[2115]<=16'd4762; ROM2[2115]<=16'd0; ROM3[2115]<=16'd23785; ROM4[2115]<=16'd57259;
ROM1[2116]<=16'd4792; ROM2[2116]<=16'd0; ROM3[2116]<=16'd23775; ROM4[2116]<=16'd57260;
ROM1[2117]<=16'd4784; ROM2[2117]<=16'd0; ROM3[2117]<=16'd23768; ROM4[2117]<=16'd57256;
ROM1[2118]<=16'd4763; ROM2[2118]<=16'd0; ROM3[2118]<=16'd23768; ROM4[2118]<=16'd57255;
ROM1[2119]<=16'd4763; ROM2[2119]<=16'd0; ROM3[2119]<=16'd23794; ROM4[2119]<=16'd57273;
ROM1[2120]<=16'd4745; ROM2[2120]<=16'd0; ROM3[2120]<=16'd23797; ROM4[2120]<=16'd57271;
ROM1[2121]<=16'd4722; ROM2[2121]<=16'd0; ROM3[2121]<=16'd23793; ROM4[2121]<=16'd57260;
ROM1[2122]<=16'd4737; ROM2[2122]<=16'd0; ROM3[2122]<=16'd23810; ROM4[2122]<=16'd57279;
ROM1[2123]<=16'd4753; ROM2[2123]<=16'd0; ROM3[2123]<=16'd23802; ROM4[2123]<=16'd57278;
ROM1[2124]<=16'd4766; ROM2[2124]<=16'd0; ROM3[2124]<=16'd23766; ROM4[2124]<=16'd57258;
ROM1[2125]<=16'd4783; ROM2[2125]<=16'd0; ROM3[2125]<=16'd23758; ROM4[2125]<=16'd57262;
ROM1[2126]<=16'd4772; ROM2[2126]<=16'd0; ROM3[2126]<=16'd23765; ROM4[2126]<=16'd57261;
ROM1[2127]<=16'd4756; ROM2[2127]<=16'd0; ROM3[2127]<=16'd23776; ROM4[2127]<=16'd57263;
ROM1[2128]<=16'd4752; ROM2[2128]<=16'd0; ROM3[2128]<=16'd23794; ROM4[2128]<=16'd57275;
ROM1[2129]<=16'd4751; ROM2[2129]<=16'd0; ROM3[2129]<=16'd23812; ROM4[2129]<=16'd57287;
ROM1[2130]<=16'd4753; ROM2[2130]<=16'd0; ROM3[2130]<=16'd23820; ROM4[2130]<=16'd57295;
ROM1[2131]<=16'd4767; ROM2[2131]<=16'd0; ROM3[2131]<=16'd23819; ROM4[2131]<=16'd57297;
ROM1[2132]<=16'd4793; ROM2[2132]<=16'd0; ROM3[2132]<=16'd23808; ROM4[2132]<=16'd57295;
ROM1[2133]<=16'd4811; ROM2[2133]<=16'd0; ROM3[2133]<=16'd23791; ROM4[2133]<=16'd57290;
ROM1[2134]<=16'd4799; ROM2[2134]<=16'd0; ROM3[2134]<=16'd23790; ROM4[2134]<=16'd57285;
ROM1[2135]<=16'd4781; ROM2[2135]<=16'd0; ROM3[2135]<=16'd23800; ROM4[2135]<=16'd57282;
ROM1[2136]<=16'd4771; ROM2[2136]<=16'd0; ROM3[2136]<=16'd23816; ROM4[2136]<=16'd57288;
ROM1[2137]<=16'd4762; ROM2[2137]<=16'd0; ROM3[2137]<=16'd23828; ROM4[2137]<=16'd57291;
ROM1[2138]<=16'd4755; ROM2[2138]<=16'd0; ROM3[2138]<=16'd23834; ROM4[2138]<=16'd57287;
ROM1[2139]<=16'd4753; ROM2[2139]<=16'd0; ROM3[2139]<=16'd23826; ROM4[2139]<=16'd57285;
ROM1[2140]<=16'd4777; ROM2[2140]<=16'd0; ROM3[2140]<=16'd23820; ROM4[2140]<=16'd57286;
ROM1[2141]<=16'd4814; ROM2[2141]<=16'd0; ROM3[2141]<=16'd23820; ROM4[2141]<=16'd57296;
ROM1[2142]<=16'd4807; ROM2[2142]<=16'd0; ROM3[2142]<=16'd23811; ROM4[2142]<=16'd57290;
ROM1[2143]<=16'd4782; ROM2[2143]<=16'd0; ROM3[2143]<=16'd23809; ROM4[2143]<=16'd57283;
ROM1[2144]<=16'd4764; ROM2[2144]<=16'd0; ROM3[2144]<=16'd23818; ROM4[2144]<=16'd57282;
ROM1[2145]<=16'd4747; ROM2[2145]<=16'd0; ROM3[2145]<=16'd23817; ROM4[2145]<=16'd57275;
ROM1[2146]<=16'd4743; ROM2[2146]<=16'd0; ROM3[2146]<=16'd23824; ROM4[2146]<=16'd57282;
ROM1[2147]<=16'd4753; ROM2[2147]<=16'd0; ROM3[2147]<=16'd23828; ROM4[2147]<=16'd57286;
ROM1[2148]<=16'd4760; ROM2[2148]<=16'd0; ROM3[2148]<=16'd23804; ROM4[2148]<=16'd57274;
ROM1[2149]<=16'd4790; ROM2[2149]<=16'd0; ROM3[2149]<=16'd23792; ROM4[2149]<=16'd57274;
ROM1[2150]<=16'd4813; ROM2[2150]<=16'd0; ROM3[2150]<=16'd23800; ROM4[2150]<=16'd57286;
ROM1[2151]<=16'd4800; ROM2[2151]<=16'd0; ROM3[2151]<=16'd23808; ROM4[2151]<=16'd57288;
ROM1[2152]<=16'd4796; ROM2[2152]<=16'd0; ROM3[2152]<=16'd23826; ROM4[2152]<=16'd57298;
ROM1[2153]<=16'd4776; ROM2[2153]<=16'd0; ROM3[2153]<=16'd23823; ROM4[2153]<=16'd57287;
ROM1[2154]<=16'd4748; ROM2[2154]<=16'd0; ROM3[2154]<=16'd23825; ROM4[2154]<=16'd57283;
ROM1[2155]<=16'd4757; ROM2[2155]<=16'd0; ROM3[2155]<=16'd23848; ROM4[2155]<=16'd57303;
ROM1[2156]<=16'd4768; ROM2[2156]<=16'd0; ROM3[2156]<=16'd23842; ROM4[2156]<=16'd57301;
ROM1[2157]<=16'd4796; ROM2[2157]<=16'd0; ROM3[2157]<=16'd23825; ROM4[2157]<=16'd57296;
ROM1[2158]<=16'd4829; ROM2[2158]<=16'd0; ROM3[2158]<=16'd23817; ROM4[2158]<=16'd57302;
ROM1[2159]<=16'd4809; ROM2[2159]<=16'd0; ROM3[2159]<=16'd23803; ROM4[2159]<=16'd57287;
ROM1[2160]<=16'd4780; ROM2[2160]<=16'd0; ROM3[2160]<=16'd23803; ROM4[2160]<=16'd57281;
ROM1[2161]<=16'd4779; ROM2[2161]<=16'd0; ROM3[2161]<=16'd23828; ROM4[2161]<=16'd57297;
ROM1[2162]<=16'd4759; ROM2[2162]<=16'd0; ROM3[2162]<=16'd23822; ROM4[2162]<=16'd57289;
ROM1[2163]<=16'd4724; ROM2[2163]<=16'd0; ROM3[2163]<=16'd23800; ROM4[2163]<=16'd57265;
ROM1[2164]<=16'd4727; ROM2[2164]<=16'd0; ROM3[2164]<=16'd23800; ROM4[2164]<=16'd57263;
ROM1[2165]<=16'd4750; ROM2[2165]<=16'd0; ROM3[2165]<=16'd23788; ROM4[2165]<=16'd57262;
ROM1[2166]<=16'd4778; ROM2[2166]<=16'd0; ROM3[2166]<=16'd23774; ROM4[2166]<=16'd57257;
ROM1[2167]<=16'd4788; ROM2[2167]<=16'd0; ROM3[2167]<=16'd23780; ROM4[2167]<=16'd57263;
ROM1[2168]<=16'd4779; ROM2[2168]<=16'd0; ROM3[2168]<=16'd23786; ROM4[2168]<=16'd57269;
ROM1[2169]<=16'd4763; ROM2[2169]<=16'd0; ROM3[2169]<=16'd23793; ROM4[2169]<=16'd57269;
ROM1[2170]<=16'd4752; ROM2[2170]<=16'd0; ROM3[2170]<=16'd23801; ROM4[2170]<=16'd57270;
ROM1[2171]<=16'd4754; ROM2[2171]<=16'd0; ROM3[2171]<=16'd23817; ROM4[2171]<=16'd57285;
ROM1[2172]<=16'd4758; ROM2[2172]<=16'd0; ROM3[2172]<=16'd23820; ROM4[2172]<=16'd57290;
ROM1[2173]<=16'd4768; ROM2[2173]<=16'd0; ROM3[2173]<=16'd23809; ROM4[2173]<=16'd57281;
ROM1[2174]<=16'd4804; ROM2[2174]<=16'd0; ROM3[2174]<=16'd23799; ROM4[2174]<=16'd57284;
ROM1[2175]<=16'd4825; ROM2[2175]<=16'd0; ROM3[2175]<=16'd23796; ROM4[2175]<=16'd57290;
ROM1[2176]<=16'd4798; ROM2[2176]<=16'd0; ROM3[2176]<=16'd23786; ROM4[2176]<=16'd57280;
ROM1[2177]<=16'd4777; ROM2[2177]<=16'd0; ROM3[2177]<=16'd23793; ROM4[2177]<=16'd57283;
ROM1[2178]<=16'd4779; ROM2[2178]<=16'd0; ROM3[2178]<=16'd23814; ROM4[2178]<=16'd57298;
ROM1[2179]<=16'd4759; ROM2[2179]<=16'd0; ROM3[2179]<=16'd23816; ROM4[2179]<=16'd57291;
ROM1[2180]<=16'd4761; ROM2[2180]<=16'd0; ROM3[2180]<=16'd23824; ROM4[2180]<=16'd57298;
ROM1[2181]<=16'd4790; ROM2[2181]<=16'd0; ROM3[2181]<=16'd23828; ROM4[2181]<=16'd57307;
ROM1[2182]<=16'd4799; ROM2[2182]<=16'd0; ROM3[2182]<=16'd23797; ROM4[2182]<=16'd57285;
ROM1[2183]<=16'd4812; ROM2[2183]<=16'd0; ROM3[2183]<=16'd23781; ROM4[2183]<=16'd57276;
ROM1[2184]<=16'd4805; ROM2[2184]<=16'd0; ROM3[2184]<=16'd23785; ROM4[2184]<=16'd57278;
ROM1[2185]<=16'd4782; ROM2[2185]<=16'd0; ROM3[2185]<=16'd23785; ROM4[2185]<=16'd57275;
ROM1[2186]<=16'd4771; ROM2[2186]<=16'd0; ROM3[2186]<=16'd23795; ROM4[2186]<=16'd57280;
ROM1[2187]<=16'd4770; ROM2[2187]<=16'd0; ROM3[2187]<=16'd23810; ROM4[2187]<=16'd57289;
ROM1[2188]<=16'd4764; ROM2[2188]<=16'd0; ROM3[2188]<=16'd23818; ROM4[2188]<=16'd57292;
ROM1[2189]<=16'd4758; ROM2[2189]<=16'd0; ROM3[2189]<=16'd23805; ROM4[2189]<=16'd57279;
ROM1[2190]<=16'd4776; ROM2[2190]<=16'd0; ROM3[2190]<=16'd23789; ROM4[2190]<=16'd57271;
ROM1[2191]<=16'd4805; ROM2[2191]<=16'd0; ROM3[2191]<=16'd23777; ROM4[2191]<=16'd57272;
ROM1[2192]<=16'd4810; ROM2[2192]<=16'd0; ROM3[2192]<=16'd23772; ROM4[2192]<=16'd57271;
ROM1[2193]<=16'd4795; ROM2[2193]<=16'd0; ROM3[2193]<=16'd23780; ROM4[2193]<=16'd57279;
ROM1[2194]<=16'd4773; ROM2[2194]<=16'd0; ROM3[2194]<=16'd23790; ROM4[2194]<=16'd57280;
ROM1[2195]<=16'd4755; ROM2[2195]<=16'd0; ROM3[2195]<=16'd23793; ROM4[2195]<=16'd57272;
ROM1[2196]<=16'd4742; ROM2[2196]<=16'd0; ROM3[2196]<=16'd23798; ROM4[2196]<=16'd57269;
ROM1[2197]<=16'd4744; ROM2[2197]<=16'd0; ROM3[2197]<=16'd23801; ROM4[2197]<=16'd57268;
ROM1[2198]<=16'd4764; ROM2[2198]<=16'd0; ROM3[2198]<=16'd23802; ROM4[2198]<=16'd57272;
ROM1[2199]<=16'd4797; ROM2[2199]<=16'd0; ROM3[2199]<=16'd23787; ROM4[2199]<=16'd57272;
ROM1[2200]<=16'd4810; ROM2[2200]<=16'd0; ROM3[2200]<=16'd23781; ROM4[2200]<=16'd57269;
ROM1[2201]<=16'd4793; ROM2[2201]<=16'd0; ROM3[2201]<=16'd23786; ROM4[2201]<=16'd57266;
ROM1[2202]<=16'd4779; ROM2[2202]<=16'd0; ROM3[2202]<=16'd23795; ROM4[2202]<=16'd57272;
ROM1[2203]<=16'd4779; ROM2[2203]<=16'd0; ROM3[2203]<=16'd23812; ROM4[2203]<=16'd57283;
ROM1[2204]<=16'd4755; ROM2[2204]<=16'd0; ROM3[2204]<=16'd23809; ROM4[2204]<=16'd57277;
ROM1[2205]<=16'd4738; ROM2[2205]<=16'd0; ROM3[2205]<=16'd23801; ROM4[2205]<=16'd57267;
ROM1[2206]<=16'd4752; ROM2[2206]<=16'd0; ROM3[2206]<=16'd23793; ROM4[2206]<=16'd57264;
ROM1[2207]<=16'd4778; ROM2[2207]<=16'd0; ROM3[2207]<=16'd23775; ROM4[2207]<=16'd57261;
ROM1[2208]<=16'd4794; ROM2[2208]<=16'd0; ROM3[2208]<=16'd23766; ROM4[2208]<=16'd57255;
ROM1[2209]<=16'd4789; ROM2[2209]<=16'd0; ROM3[2209]<=16'd23769; ROM4[2209]<=16'd57259;
ROM1[2210]<=16'd4761; ROM2[2210]<=16'd0; ROM3[2210]<=16'd23766; ROM4[2210]<=16'd57254;
ROM1[2211]<=16'd4741; ROM2[2211]<=16'd0; ROM3[2211]<=16'd23776; ROM4[2211]<=16'd57257;
ROM1[2212]<=16'd4733; ROM2[2212]<=16'd0; ROM3[2212]<=16'd23786; ROM4[2212]<=16'd57264;
ROM1[2213]<=16'd4709; ROM2[2213]<=16'd0; ROM3[2213]<=16'd23770; ROM4[2213]<=16'd57246;
ROM1[2214]<=16'd4706; ROM2[2214]<=16'd0; ROM3[2214]<=16'd23761; ROM4[2214]<=16'd57234;
ROM1[2215]<=16'd4736; ROM2[2215]<=16'd0; ROM3[2215]<=16'd23757; ROM4[2215]<=16'd57237;
ROM1[2216]<=16'd4774; ROM2[2216]<=16'd0; ROM3[2216]<=16'd23760; ROM4[2216]<=16'd57252;
ROM1[2217]<=16'd4793; ROM2[2217]<=16'd0; ROM3[2217]<=16'd23780; ROM4[2217]<=16'd57274;
ROM1[2218]<=16'd4790; ROM2[2218]<=16'd0; ROM3[2218]<=16'd23800; ROM4[2218]<=16'd57287;
ROM1[2219]<=16'd4771; ROM2[2219]<=16'd0; ROM3[2219]<=16'd23811; ROM4[2219]<=16'd57287;
ROM1[2220]<=16'd4744; ROM2[2220]<=16'd0; ROM3[2220]<=16'd23804; ROM4[2220]<=16'd57271;
ROM1[2221]<=16'd4723; ROM2[2221]<=16'd0; ROM3[2221]<=16'd23803; ROM4[2221]<=16'd57263;
ROM1[2222]<=16'd4728; ROM2[2222]<=16'd0; ROM3[2222]<=16'd23805; ROM4[2222]<=16'd57268;
ROM1[2223]<=16'd4746; ROM2[2223]<=16'd0; ROM3[2223]<=16'd23792; ROM4[2223]<=16'd57265;
ROM1[2224]<=16'd4776; ROM2[2224]<=16'd0; ROM3[2224]<=16'd23775; ROM4[2224]<=16'd57266;
ROM1[2225]<=16'd4797; ROM2[2225]<=16'd0; ROM3[2225]<=16'd23774; ROM4[2225]<=16'd57273;
ROM1[2226]<=16'd4788; ROM2[2226]<=16'd0; ROM3[2226]<=16'd23782; ROM4[2226]<=16'd57278;
ROM1[2227]<=16'd4767; ROM2[2227]<=16'd0; ROM3[2227]<=16'd23785; ROM4[2227]<=16'd57279;
ROM1[2228]<=16'd4760; ROM2[2228]<=16'd0; ROM3[2228]<=16'd23790; ROM4[2228]<=16'd57281;
ROM1[2229]<=16'd4747; ROM2[2229]<=16'd0; ROM3[2229]<=16'd23794; ROM4[2229]<=16'd57278;
ROM1[2230]<=16'd4734; ROM2[2230]<=16'd0; ROM3[2230]<=16'd23789; ROM4[2230]<=16'd57269;
ROM1[2231]<=16'd4742; ROM2[2231]<=16'd0; ROM3[2231]<=16'd23782; ROM4[2231]<=16'd57263;
ROM1[2232]<=16'd4767; ROM2[2232]<=16'd0; ROM3[2232]<=16'd23775; ROM4[2232]<=16'd57261;
ROM1[2233]<=16'd4790; ROM2[2233]<=16'd0; ROM3[2233]<=16'd23768; ROM4[2233]<=16'd57263;
ROM1[2234]<=16'd4784; ROM2[2234]<=16'd0; ROM3[2234]<=16'd23771; ROM4[2234]<=16'd57258;
ROM1[2235]<=16'd4754; ROM2[2235]<=16'd0; ROM3[2235]<=16'd23764; ROM4[2235]<=16'd57244;
ROM1[2236]<=16'd4739; ROM2[2236]<=16'd0; ROM3[2236]<=16'd23766; ROM4[2236]<=16'd57241;
ROM1[2237]<=16'd4723; ROM2[2237]<=16'd0; ROM3[2237]<=16'd23767; ROM4[2237]<=16'd57237;
ROM1[2238]<=16'd4708; ROM2[2238]<=16'd0; ROM3[2238]<=16'd23764; ROM4[2238]<=16'd57235;
ROM1[2239]<=16'd4721; ROM2[2239]<=16'd0; ROM3[2239]<=16'd23768; ROM4[2239]<=16'd57241;
ROM1[2240]<=16'd4742; ROM2[2240]<=16'd0; ROM3[2240]<=16'd23758; ROM4[2240]<=16'd57241;
ROM1[2241]<=16'd4772; ROM2[2241]<=16'd0; ROM3[2241]<=16'd23744; ROM4[2241]<=16'd57240;
ROM1[2242]<=16'd4793; ROM2[2242]<=16'd0; ROM3[2242]<=16'd23756; ROM4[2242]<=16'd57256;
ROM1[2243]<=16'd4784; ROM2[2243]<=16'd0; ROM3[2243]<=16'd23764; ROM4[2243]<=16'd57265;
ROM1[2244]<=16'd4754; ROM2[2244]<=16'd0; ROM3[2244]<=16'd23760; ROM4[2244]<=16'd57253;
ROM1[2245]<=16'd4738; ROM2[2245]<=16'd0; ROM3[2245]<=16'd23767; ROM4[2245]<=16'd57251;
ROM1[2246]<=16'd4714; ROM2[2246]<=16'd0; ROM3[2246]<=16'd23760; ROM4[2246]<=16'd57241;
ROM1[2247]<=16'd4708; ROM2[2247]<=16'd0; ROM3[2247]<=16'd23757; ROM4[2247]<=16'd57236;
ROM1[2248]<=16'd4739; ROM2[2248]<=16'd0; ROM3[2248]<=16'd23762; ROM4[2248]<=16'd57248;
ROM1[2249]<=16'd4768; ROM2[2249]<=16'd0; ROM3[2249]<=16'd23742; ROM4[2249]<=16'd57244;
ROM1[2250]<=16'd4765; ROM2[2250]<=16'd0; ROM3[2250]<=16'd23722; ROM4[2250]<=16'd57230;
ROM1[2251]<=16'd4757; ROM2[2251]<=16'd0; ROM3[2251]<=16'd23733; ROM4[2251]<=16'd57234;
ROM1[2252]<=16'd4759; ROM2[2252]<=16'd0; ROM3[2252]<=16'd23759; ROM4[2252]<=16'd57253;
ROM1[2253]<=16'd4740; ROM2[2253]<=16'd0; ROM3[2253]<=16'd23761; ROM4[2253]<=16'd57247;
ROM1[2254]<=16'd4712; ROM2[2254]<=16'd0; ROM3[2254]<=16'd23756; ROM4[2254]<=16'd57237;
ROM1[2255]<=16'd4708; ROM2[2255]<=16'd0; ROM3[2255]<=16'd23761; ROM4[2255]<=16'd57238;
ROM1[2256]<=16'd4719; ROM2[2256]<=16'd0; ROM3[2256]<=16'd23751; ROM4[2256]<=16'd57231;
ROM1[2257]<=16'd4750; ROM2[2257]<=16'd0; ROM3[2257]<=16'd23740; ROM4[2257]<=16'd57232;
ROM1[2258]<=16'd4775; ROM2[2258]<=16'd0; ROM3[2258]<=16'd23736; ROM4[2258]<=16'd57240;
ROM1[2259]<=16'd4768; ROM2[2259]<=16'd0; ROM3[2259]<=16'd23740; ROM4[2259]<=16'd57243;
ROM1[2260]<=16'd4741; ROM2[2260]<=16'd0; ROM3[2260]<=16'd23743; ROM4[2260]<=16'd57235;
ROM1[2261]<=16'd4717; ROM2[2261]<=16'd0; ROM3[2261]<=16'd23742; ROM4[2261]<=16'd57228;
ROM1[2262]<=16'd4712; ROM2[2262]<=16'd0; ROM3[2262]<=16'd23756; ROM4[2262]<=16'd57235;
ROM1[2263]<=16'd4714; ROM2[2263]<=16'd0; ROM3[2263]<=16'd23767; ROM4[2263]<=16'd57241;
ROM1[2264]<=16'd4733; ROM2[2264]<=16'd0; ROM3[2264]<=16'd23776; ROM4[2264]<=16'd57256;
ROM1[2265]<=16'd4761; ROM2[2265]<=16'd0; ROM3[2265]<=16'd23772; ROM4[2265]<=16'd57263;
ROM1[2266]<=16'd4769; ROM2[2266]<=16'd0; ROM3[2266]<=16'd23740; ROM4[2266]<=16'd57240;
ROM1[2267]<=16'd4754; ROM2[2267]<=16'd0; ROM3[2267]<=16'd23720; ROM4[2267]<=16'd57222;
ROM1[2268]<=16'd4732; ROM2[2268]<=16'd0; ROM3[2268]<=16'd23717; ROM4[2268]<=16'd57216;
ROM1[2269]<=16'd4717; ROM2[2269]<=16'd0; ROM3[2269]<=16'd23733; ROM4[2269]<=16'd57221;
ROM1[2270]<=16'd4714; ROM2[2270]<=16'd0; ROM3[2270]<=16'd23755; ROM4[2270]<=16'd57233;
ROM1[2271]<=16'd4705; ROM2[2271]<=16'd0; ROM3[2271]<=16'd23771; ROM4[2271]<=16'd57242;
ROM1[2272]<=16'd4701; ROM2[2272]<=16'd0; ROM3[2272]<=16'd23763; ROM4[2272]<=16'd57236;
ROM1[2273]<=16'd4709; ROM2[2273]<=16'd0; ROM3[2273]<=16'd23735; ROM4[2273]<=16'd57215;
ROM1[2274]<=16'd4743; ROM2[2274]<=16'd0; ROM3[2274]<=16'd23721; ROM4[2274]<=16'd57213;
ROM1[2275]<=16'd4747; ROM2[2275]<=16'd0; ROM3[2275]<=16'd23705; ROM4[2275]<=16'd57207;
ROM1[2276]<=16'd4728; ROM2[2276]<=16'd0; ROM3[2276]<=16'd23711; ROM4[2276]<=16'd57206;
ROM1[2277]<=16'd4728; ROM2[2277]<=16'd0; ROM3[2277]<=16'd23745; ROM4[2277]<=16'd57229;
ROM1[2278]<=16'd4727; ROM2[2278]<=16'd0; ROM3[2278]<=16'd23767; ROM4[2278]<=16'd57246;
ROM1[2279]<=16'd4730; ROM2[2279]<=16'd0; ROM3[2279]<=16'd23787; ROM4[2279]<=16'd57262;
ROM1[2280]<=16'd4728; ROM2[2280]<=16'd0; ROM3[2280]<=16'd23787; ROM4[2280]<=16'd57262;
ROM1[2281]<=16'd4723; ROM2[2281]<=16'd0; ROM3[2281]<=16'd23765; ROM4[2281]<=16'd57246;
ROM1[2282]<=16'd4732; ROM2[2282]<=16'd0; ROM3[2282]<=16'd23733; ROM4[2282]<=16'd57223;
ROM1[2283]<=16'd4740; ROM2[2283]<=16'd0; ROM3[2283]<=16'd23715; ROM4[2283]<=16'd57211;
ROM1[2284]<=16'd4734; ROM2[2284]<=16'd0; ROM3[2284]<=16'd23722; ROM4[2284]<=16'd57214;
ROM1[2285]<=16'd4724; ROM2[2285]<=16'd0; ROM3[2285]<=16'd23737; ROM4[2285]<=16'd57218;
ROM1[2286]<=16'd4715; ROM2[2286]<=16'd0; ROM3[2286]<=16'd23752; ROM4[2286]<=16'd57224;
ROM1[2287]<=16'd4695; ROM2[2287]<=16'd0; ROM3[2287]<=16'd23757; ROM4[2287]<=16'd57221;
ROM1[2288]<=16'd4678; ROM2[2288]<=16'd0; ROM3[2288]<=16'd23755; ROM4[2288]<=16'd57216;
ROM1[2289]<=16'd4680; ROM2[2289]<=16'd0; ROM3[2289]<=16'd23752; ROM4[2289]<=16'd57213;
ROM1[2290]<=16'd4716; ROM2[2290]<=16'd0; ROM3[2290]<=16'd23750; ROM4[2290]<=16'd57223;
ROM1[2291]<=16'd4763; ROM2[2291]<=16'd0; ROM3[2291]<=16'd23747; ROM4[2291]<=16'd57236;
ROM1[2292]<=16'd4754; ROM2[2292]<=16'd0; ROM3[2292]<=16'd23738; ROM4[2292]<=16'd57228;
ROM1[2293]<=16'd4730; ROM2[2293]<=16'd0; ROM3[2293]<=16'd23733; ROM4[2293]<=16'd57217;
ROM1[2294]<=16'd4711; ROM2[2294]<=16'd0; ROM3[2294]<=16'd23743; ROM4[2294]<=16'd57217;
ROM1[2295]<=16'd4693; ROM2[2295]<=16'd0; ROM3[2295]<=16'd23749; ROM4[2295]<=16'd57216;
ROM1[2296]<=16'd4691; ROM2[2296]<=16'd0; ROM3[2296]<=16'd23763; ROM4[2296]<=16'd57228;
ROM1[2297]<=16'd4702; ROM2[2297]<=16'd0; ROM3[2297]<=16'd23773; ROM4[2297]<=16'd57240;
ROM1[2298]<=16'd4721; ROM2[2298]<=16'd0; ROM3[2298]<=16'd23765; ROM4[2298]<=16'd57240;
ROM1[2299]<=16'd4748; ROM2[2299]<=16'd0; ROM3[2299]<=16'd23748; ROM4[2299]<=16'd57236;
ROM1[2300]<=16'd4751; ROM2[2300]<=16'd0; ROM3[2300]<=16'd23732; ROM4[2300]<=16'd57227;
ROM1[2301]<=16'd4742; ROM2[2301]<=16'd0; ROM3[2301]<=16'd23738; ROM4[2301]<=16'd57235;
ROM1[2302]<=16'd4738; ROM2[2302]<=16'd0; ROM3[2302]<=16'd23759; ROM4[2302]<=16'd57249;
ROM1[2303]<=16'd4723; ROM2[2303]<=16'd0; ROM3[2303]<=16'd23762; ROM4[2303]<=16'd57244;
ROM1[2304]<=16'd4711; ROM2[2304]<=16'd0; ROM3[2304]<=16'd23771; ROM4[2304]<=16'd57251;
ROM1[2305]<=16'd4717; ROM2[2305]<=16'd0; ROM3[2305]<=16'd23787; ROM4[2305]<=16'd57262;
ROM1[2306]<=16'd4719; ROM2[2306]<=16'd0; ROM3[2306]<=16'd23774; ROM4[2306]<=16'd57248;
ROM1[2307]<=16'd4745; ROM2[2307]<=16'd0; ROM3[2307]<=16'd23760; ROM4[2307]<=16'd57247;
ROM1[2308]<=16'd4775; ROM2[2308]<=16'd0; ROM3[2308]<=16'd23757; ROM4[2308]<=16'd57254;
ROM1[2309]<=16'd4768; ROM2[2309]<=16'd0; ROM3[2309]<=16'd23759; ROM4[2309]<=16'd57253;
ROM1[2310]<=16'd4760; ROM2[2310]<=16'd0; ROM3[2310]<=16'd23771; ROM4[2310]<=16'd57263;
ROM1[2311]<=16'd4742; ROM2[2311]<=16'd0; ROM3[2311]<=16'd23778; ROM4[2311]<=16'd57259;
ROM1[2312]<=16'd4726; ROM2[2312]<=16'd0; ROM3[2312]<=16'd23783; ROM4[2312]<=16'd57258;
ROM1[2313]<=16'd4728; ROM2[2313]<=16'd0; ROM3[2313]<=16'd23800; ROM4[2313]<=16'd57273;
ROM1[2314]<=16'd4736; ROM2[2314]<=16'd0; ROM3[2314]<=16'd23802; ROM4[2314]<=16'd57275;
ROM1[2315]<=16'd4756; ROM2[2315]<=16'd0; ROM3[2315]<=16'd23786; ROM4[2315]<=16'd57273;
ROM1[2316]<=16'd4774; ROM2[2316]<=16'd0; ROM3[2316]<=16'd23766; ROM4[2316]<=16'd57261;
ROM1[2317]<=16'd4760; ROM2[2317]<=16'd0; ROM3[2317]<=16'd23744; ROM4[2317]<=16'd57239;
ROM1[2318]<=16'd4722; ROM2[2318]<=16'd0; ROM3[2318]<=16'd23728; ROM4[2318]<=16'd57217;
ROM1[2319]<=16'd4710; ROM2[2319]<=16'd0; ROM3[2319]<=16'd23743; ROM4[2319]<=16'd57220;
ROM1[2320]<=16'd4729; ROM2[2320]<=16'd0; ROM3[2320]<=16'd23768; ROM4[2320]<=16'd57245;
ROM1[2321]<=16'd4698; ROM2[2321]<=16'd0; ROM3[2321]<=16'd23756; ROM4[2321]<=16'd57230;
ROM1[2322]<=16'd4680; ROM2[2322]<=16'd0; ROM3[2322]<=16'd23745; ROM4[2322]<=16'd57218;
ROM1[2323]<=16'd4696; ROM2[2323]<=16'd0; ROM3[2323]<=16'd23736; ROM4[2323]<=16'd57216;
ROM1[2324]<=16'd4725; ROM2[2324]<=16'd0; ROM3[2324]<=16'd23722; ROM4[2324]<=16'd57209;
ROM1[2325]<=16'd4755; ROM2[2325]<=16'd0; ROM3[2325]<=16'd23728; ROM4[2325]<=16'd57222;
ROM1[2326]<=16'd4752; ROM2[2326]<=16'd0; ROM3[2326]<=16'd23737; ROM4[2326]<=16'd57231;
ROM1[2327]<=16'd4734; ROM2[2327]<=16'd0; ROM3[2327]<=16'd23747; ROM4[2327]<=16'd57233;
ROM1[2328]<=16'd4717; ROM2[2328]<=16'd0; ROM3[2328]<=16'd23758; ROM4[2328]<=16'd57236;
ROM1[2329]<=16'd4702; ROM2[2329]<=16'd0; ROM3[2329]<=16'd23770; ROM4[2329]<=16'd57239;
ROM1[2330]<=16'd4697; ROM2[2330]<=16'd0; ROM3[2330]<=16'd23770; ROM4[2330]<=16'd57236;
ROM1[2331]<=16'd4712; ROM2[2331]<=16'd0; ROM3[2331]<=16'd23762; ROM4[2331]<=16'd57235;
ROM1[2332]<=16'd4738; ROM2[2332]<=16'd0; ROM3[2332]<=16'd23744; ROM4[2332]<=16'd57227;
ROM1[2333]<=16'd4756; ROM2[2333]<=16'd0; ROM3[2333]<=16'd23726; ROM4[2333]<=16'd57221;
ROM1[2334]<=16'd4756; ROM2[2334]<=16'd0; ROM3[2334]<=16'd23733; ROM4[2334]<=16'd57227;
ROM1[2335]<=16'd4725; ROM2[2335]<=16'd0; ROM3[2335]<=16'd23731; ROM4[2335]<=16'd57217;
ROM1[2336]<=16'd4705; ROM2[2336]<=16'd0; ROM3[2336]<=16'd23734; ROM4[2336]<=16'd57210;
ROM1[2337]<=16'd4695; ROM2[2337]<=16'd0; ROM3[2337]<=16'd23747; ROM4[2337]<=16'd57213;
ROM1[2338]<=16'd4694; ROM2[2338]<=16'd0; ROM3[2338]<=16'd23766; ROM4[2338]<=16'd57224;
ROM1[2339]<=16'd4716; ROM2[2339]<=16'd0; ROM3[2339]<=16'd23775; ROM4[2339]<=16'd57239;
ROM1[2340]<=16'd4721; ROM2[2340]<=16'd0; ROM3[2340]<=16'd23748; ROM4[2340]<=16'd57222;
ROM1[2341]<=16'd4749; ROM2[2341]<=16'd0; ROM3[2341]<=16'd23736; ROM4[2341]<=16'd57219;
ROM1[2342]<=16'd4759; ROM2[2342]<=16'd0; ROM3[2342]<=16'd23738; ROM4[2342]<=16'd57230;
ROM1[2343]<=16'd4741; ROM2[2343]<=16'd0; ROM3[2343]<=16'd23744; ROM4[2343]<=16'd57230;
ROM1[2344]<=16'd4736; ROM2[2344]<=16'd0; ROM3[2344]<=16'd23765; ROM4[2344]<=16'd57244;
ROM1[2345]<=16'd4729; ROM2[2345]<=16'd0; ROM3[2345]<=16'd23777; ROM4[2345]<=16'd57253;
ROM1[2346]<=16'd4711; ROM2[2346]<=16'd0; ROM3[2346]<=16'd23780; ROM4[2346]<=16'd57248;
ROM1[2347]<=16'd4718; ROM2[2347]<=16'd0; ROM3[2347]<=16'd23797; ROM4[2347]<=16'd57255;
ROM1[2348]<=16'd4743; ROM2[2348]<=16'd0; ROM3[2348]<=16'd23796; ROM4[2348]<=16'd57262;
ROM1[2349]<=16'd4763; ROM2[2349]<=16'd0; ROM3[2349]<=16'd23767; ROM4[2349]<=16'd57252;
ROM1[2350]<=16'd4764; ROM2[2350]<=16'd0; ROM3[2350]<=16'd23752; ROM4[2350]<=16'd57237;
ROM1[2351]<=16'd4750; ROM2[2351]<=16'd0; ROM3[2351]<=16'd23752; ROM4[2351]<=16'd57230;
ROM1[2352]<=16'd4732; ROM2[2352]<=16'd0; ROM3[2352]<=16'd23761; ROM4[2352]<=16'd57232;
ROM1[2353]<=16'd4725; ROM2[2353]<=16'd0; ROM3[2353]<=16'd23775; ROM4[2353]<=16'd57242;
ROM1[2354]<=16'd4711; ROM2[2354]<=16'd0; ROM3[2354]<=16'd23783; ROM4[2354]<=16'd57247;
ROM1[2355]<=16'd4699; ROM2[2355]<=16'd0; ROM3[2355]<=16'd23782; ROM4[2355]<=16'd57245;
ROM1[2356]<=16'd4717; ROM2[2356]<=16'd0; ROM3[2356]<=16'd23781; ROM4[2356]<=16'd57248;
ROM1[2357]<=16'd4755; ROM2[2357]<=16'd0; ROM3[2357]<=16'd23774; ROM4[2357]<=16'd57252;
ROM1[2358]<=16'd4788; ROM2[2358]<=16'd0; ROM3[2358]<=16'd23772; ROM4[2358]<=16'd57260;
ROM1[2359]<=16'd4794; ROM2[2359]<=16'd0; ROM3[2359]<=16'd23779; ROM4[2359]<=16'd57273;
ROM1[2360]<=16'd4766; ROM2[2360]<=16'd0; ROM3[2360]<=16'd23778; ROM4[2360]<=16'd57262;
ROM1[2361]<=16'd4724; ROM2[2361]<=16'd0; ROM3[2361]<=16'd23757; ROM4[2361]<=16'd57236;
ROM1[2362]<=16'd4701; ROM2[2362]<=16'd0; ROM3[2362]<=16'd23744; ROM4[2362]<=16'd57225;
ROM1[2363]<=16'd4696; ROM2[2363]<=16'd0; ROM3[2363]<=16'd23754; ROM4[2363]<=16'd57233;
ROM1[2364]<=16'd4713; ROM2[2364]<=16'd0; ROM3[2364]<=16'd23766; ROM4[2364]<=16'd57245;
ROM1[2365]<=16'd4737; ROM2[2365]<=16'd0; ROM3[2365]<=16'd23754; ROM4[2365]<=16'd57242;
ROM1[2366]<=16'd4759; ROM2[2366]<=16'd0; ROM3[2366]<=16'd23740; ROM4[2366]<=16'd57237;
ROM1[2367]<=16'd4761; ROM2[2367]<=16'd0; ROM3[2367]<=16'd23733; ROM4[2367]<=16'd57232;
ROM1[2368]<=16'd4748; ROM2[2368]<=16'd0; ROM3[2368]<=16'd23746; ROM4[2368]<=16'd57236;
ROM1[2369]<=16'd4753; ROM2[2369]<=16'd0; ROM3[2369]<=16'd23784; ROM4[2369]<=16'd57261;
ROM1[2370]<=16'd4747; ROM2[2370]<=16'd0; ROM3[2370]<=16'd23797; ROM4[2370]<=16'd57270;
ROM1[2371]<=16'd4720; ROM2[2371]<=16'd0; ROM3[2371]<=16'd23790; ROM4[2371]<=16'd57259;
ROM1[2372]<=16'd4718; ROM2[2372]<=16'd0; ROM3[2372]<=16'd23784; ROM4[2372]<=16'd57254;
ROM1[2373]<=16'd4757; ROM2[2373]<=16'd0; ROM3[2373]<=16'd23797; ROM4[2373]<=16'd57274;
ROM1[2374]<=16'd4802; ROM2[2374]<=16'd0; ROM3[2374]<=16'd23804; ROM4[2374]<=16'd57289;
ROM1[2375]<=16'd4801; ROM2[2375]<=16'd0; ROM3[2375]<=16'd23792; ROM4[2375]<=16'd57277;
ROM1[2376]<=16'd4760; ROM2[2376]<=16'd0; ROM3[2376]<=16'd23767; ROM4[2376]<=16'd57251;
ROM1[2377]<=16'd4730; ROM2[2377]<=16'd0; ROM3[2377]<=16'd23760; ROM4[2377]<=16'd57244;
ROM1[2378]<=16'd4726; ROM2[2378]<=16'd0; ROM3[2378]<=16'd23778; ROM4[2378]<=16'd57255;
ROM1[2379]<=16'd4726; ROM2[2379]<=16'd0; ROM3[2379]<=16'd23800; ROM4[2379]<=16'd57269;
ROM1[2380]<=16'd4742; ROM2[2380]<=16'd0; ROM3[2380]<=16'd23825; ROM4[2380]<=16'd57294;
ROM1[2381]<=16'd4747; ROM2[2381]<=16'd0; ROM3[2381]<=16'd23812; ROM4[2381]<=16'd57285;
ROM1[2382]<=16'd4758; ROM2[2382]<=16'd0; ROM3[2382]<=16'd23783; ROM4[2382]<=16'd57265;
ROM1[2383]<=16'd4781; ROM2[2383]<=16'd0; ROM3[2383]<=16'd23773; ROM4[2383]<=16'd57270;
ROM1[2384]<=16'd4777; ROM2[2384]<=16'd0; ROM3[2384]<=16'd23771; ROM4[2384]<=16'd57269;
ROM1[2385]<=16'd4761; ROM2[2385]<=16'd0; ROM3[2385]<=16'd23777; ROM4[2385]<=16'd57265;
ROM1[2386]<=16'd4755; ROM2[2386]<=16'd0; ROM3[2386]<=16'd23790; ROM4[2386]<=16'd57269;
ROM1[2387]<=16'd4745; ROM2[2387]<=16'd0; ROM3[2387]<=16'd23797; ROM4[2387]<=16'd57270;
ROM1[2388]<=16'd4727; ROM2[2388]<=16'd0; ROM3[2388]<=16'd23794; ROM4[2388]<=16'd57263;
ROM1[2389]<=16'd4734; ROM2[2389]<=16'd0; ROM3[2389]<=16'd23792; ROM4[2389]<=16'd57262;
ROM1[2390]<=16'd4756; ROM2[2390]<=16'd0; ROM3[2390]<=16'd23774; ROM4[2390]<=16'd57255;
ROM1[2391]<=16'd4784; ROM2[2391]<=16'd0; ROM3[2391]<=16'd23758; ROM4[2391]<=16'd57249;
ROM1[2392]<=16'd4791; ROM2[2392]<=16'd0; ROM3[2392]<=16'd23772; ROM4[2392]<=16'd57260;
ROM1[2393]<=16'd4779; ROM2[2393]<=16'd0; ROM3[2393]<=16'd23788; ROM4[2393]<=16'd57268;
ROM1[2394]<=16'd4749; ROM2[2394]<=16'd0; ROM3[2394]<=16'd23785; ROM4[2394]<=16'd57260;
ROM1[2395]<=16'd4721; ROM2[2395]<=16'd0; ROM3[2395]<=16'd23779; ROM4[2395]<=16'd57251;
ROM1[2396]<=16'd4704; ROM2[2396]<=16'd0; ROM3[2396]<=16'd23777; ROM4[2396]<=16'd57246;
ROM1[2397]<=16'd4702; ROM2[2397]<=16'd0; ROM3[2397]<=16'd23770; ROM4[2397]<=16'd57238;
ROM1[2398]<=16'd4723; ROM2[2398]<=16'd0; ROM3[2398]<=16'd23763; ROM4[2398]<=16'd57236;
ROM1[2399]<=16'd4758; ROM2[2399]<=16'd0; ROM3[2399]<=16'd23753; ROM4[2399]<=16'd57240;
ROM1[2400]<=16'd4770; ROM2[2400]<=16'd0; ROM3[2400]<=16'd23751; ROM4[2400]<=16'd57240;
ROM1[2401]<=16'd4763; ROM2[2401]<=16'd0; ROM3[2401]<=16'd23762; ROM4[2401]<=16'd57245;
ROM1[2402]<=16'd4744; ROM2[2402]<=16'd0; ROM3[2402]<=16'd23773; ROM4[2402]<=16'd57247;
ROM1[2403]<=16'd4732; ROM2[2403]<=16'd0; ROM3[2403]<=16'd23785; ROM4[2403]<=16'd57250;
ROM1[2404]<=16'd4732; ROM2[2404]<=16'd0; ROM3[2404]<=16'd23802; ROM4[2404]<=16'd57264;
ROM1[2405]<=16'd4724; ROM2[2405]<=16'd0; ROM3[2405]<=16'd23800; ROM4[2405]<=16'd57258;
ROM1[2406]<=16'd4733; ROM2[2406]<=16'd0; ROM3[2406]<=16'd23787; ROM4[2406]<=16'd57253;
ROM1[2407]<=16'd4762; ROM2[2407]<=16'd0; ROM3[2407]<=16'd23772; ROM4[2407]<=16'd57251;
ROM1[2408]<=16'd4773; ROM2[2408]<=16'd0; ROM3[2408]<=16'd23754; ROM4[2408]<=16'd57239;
ROM1[2409]<=16'd4768; ROM2[2409]<=16'd0; ROM3[2409]<=16'd23769; ROM4[2409]<=16'd57247;
ROM1[2410]<=16'd4756; ROM2[2410]<=16'd0; ROM3[2410]<=16'd23785; ROM4[2410]<=16'd57256;
ROM1[2411]<=16'd4739; ROM2[2411]<=16'd0; ROM3[2411]<=16'd23789; ROM4[2411]<=16'd57255;
ROM1[2412]<=16'd4729; ROM2[2412]<=16'd0; ROM3[2412]<=16'd23791; ROM4[2412]<=16'd57257;
ROM1[2413]<=16'd4721; ROM2[2413]<=16'd0; ROM3[2413]<=16'd23792; ROM4[2413]<=16'd57258;
ROM1[2414]<=16'd4729; ROM2[2414]<=16'd0; ROM3[2414]<=16'd23790; ROM4[2414]<=16'd57261;
ROM1[2415]<=16'd4752; ROM2[2415]<=16'd0; ROM3[2415]<=16'd23780; ROM4[2415]<=16'd57262;
ROM1[2416]<=16'd4783; ROM2[2416]<=16'd0; ROM3[2416]<=16'd23772; ROM4[2416]<=16'd57262;
ROM1[2417]<=16'd4800; ROM2[2417]<=16'd0; ROM3[2417]<=16'd23781; ROM4[2417]<=16'd57274;
ROM1[2418]<=16'd4787; ROM2[2418]<=16'd0; ROM3[2418]<=16'd23791; ROM4[2418]<=16'd57277;
ROM1[2419]<=16'd4758; ROM2[2419]<=16'd0; ROM3[2419]<=16'd23792; ROM4[2419]<=16'd57266;
ROM1[2420]<=16'd4743; ROM2[2420]<=16'd0; ROM3[2420]<=16'd23792; ROM4[2420]<=16'd57263;
ROM1[2421]<=16'd4714; ROM2[2421]<=16'd0; ROM3[2421]<=16'd23782; ROM4[2421]<=16'd57251;
ROM1[2422]<=16'd4718; ROM2[2422]<=16'd0; ROM3[2422]<=16'd23785; ROM4[2422]<=16'd57251;
ROM1[2423]<=16'd4755; ROM2[2423]<=16'd0; ROM3[2423]<=16'd23790; ROM4[2423]<=16'd57263;
ROM1[2424]<=16'd4783; ROM2[2424]<=16'd0; ROM3[2424]<=16'd23784; ROM4[2424]<=16'd57264;
ROM1[2425]<=16'd4796; ROM2[2425]<=16'd0; ROM3[2425]<=16'd23786; ROM4[2425]<=16'd57272;
ROM1[2426]<=16'd4795; ROM2[2426]<=16'd0; ROM3[2426]<=16'd23802; ROM4[2426]<=16'd57289;
ROM1[2427]<=16'd4784; ROM2[2427]<=16'd0; ROM3[2427]<=16'd23819; ROM4[2427]<=16'd57294;
ROM1[2428]<=16'd4761; ROM2[2428]<=16'd0; ROM3[2428]<=16'd23811; ROM4[2428]<=16'd57281;
ROM1[2429]<=16'd4747; ROM2[2429]<=16'd0; ROM3[2429]<=16'd23816; ROM4[2429]<=16'd57282;
ROM1[2430]<=16'd4744; ROM2[2430]<=16'd0; ROM3[2430]<=16'd23820; ROM4[2430]<=16'd57285;
ROM1[2431]<=16'd4745; ROM2[2431]<=16'd0; ROM3[2431]<=16'd23796; ROM4[2431]<=16'd57272;
ROM1[2432]<=16'd4783; ROM2[2432]<=16'd0; ROM3[2432]<=16'd23787; ROM4[2432]<=16'd57279;
ROM1[2433]<=16'd4812; ROM2[2433]<=16'd0; ROM3[2433]<=16'd23785; ROM4[2433]<=16'd57287;
ROM1[2434]<=16'd4793; ROM2[2434]<=16'd0; ROM3[2434]<=16'd23774; ROM4[2434]<=16'd57272;
ROM1[2435]<=16'd4768; ROM2[2435]<=16'd0; ROM3[2435]<=16'd23774; ROM4[2435]<=16'd57263;
ROM1[2436]<=16'd4757; ROM2[2436]<=16'd0; ROM3[2436]<=16'd23785; ROM4[2436]<=16'd57267;
ROM1[2437]<=16'd4742; ROM2[2437]<=16'd0; ROM3[2437]<=16'd23789; ROM4[2437]<=16'd57266;
ROM1[2438]<=16'd4732; ROM2[2438]<=16'd0; ROM3[2438]<=16'd23790; ROM4[2438]<=16'd57265;
ROM1[2439]<=16'd4749; ROM2[2439]<=16'd0; ROM3[2439]<=16'd23800; ROM4[2439]<=16'd57274;
ROM1[2440]<=16'd4771; ROM2[2440]<=16'd0; ROM3[2440]<=16'd23792; ROM4[2440]<=16'd57275;
ROM1[2441]<=16'd4793; ROM2[2441]<=16'd0; ROM3[2441]<=16'd23776; ROM4[2441]<=16'd57268;
ROM1[2442]<=16'd4789; ROM2[2442]<=16'd0; ROM3[2442]<=16'd23776; ROM4[2442]<=16'd57266;
ROM1[2443]<=16'd4772; ROM2[2443]<=16'd0; ROM3[2443]<=16'd23784; ROM4[2443]<=16'd57272;
ROM1[2444]<=16'd4751; ROM2[2444]<=16'd0; ROM3[2444]<=16'd23790; ROM4[2444]<=16'd57271;
ROM1[2445]<=16'd4729; ROM2[2445]<=16'd0; ROM3[2445]<=16'd23785; ROM4[2445]<=16'd57263;
ROM1[2446]<=16'd4716; ROM2[2446]<=16'd0; ROM3[2446]<=16'd23782; ROM4[2446]<=16'd57258;
ROM1[2447]<=16'd4718; ROM2[2447]<=16'd0; ROM3[2447]<=16'd23780; ROM4[2447]<=16'd57257;
ROM1[2448]<=16'd4737; ROM2[2448]<=16'd0; ROM3[2448]<=16'd23771; ROM4[2448]<=16'd57257;
ROM1[2449]<=16'd4773; ROM2[2449]<=16'd0; ROM3[2449]<=16'd23759; ROM4[2449]<=16'd57263;
ROM1[2450]<=16'd4779; ROM2[2450]<=16'd0; ROM3[2450]<=16'd23756; ROM4[2450]<=16'd57262;
ROM1[2451]<=16'd4765; ROM2[2451]<=16'd0; ROM3[2451]<=16'd23763; ROM4[2451]<=16'd57262;
ROM1[2452]<=16'd4755; ROM2[2452]<=16'd0; ROM3[2452]<=16'd23773; ROM4[2452]<=16'd57267;
ROM1[2453]<=16'd4740; ROM2[2453]<=16'd0; ROM3[2453]<=16'd23776; ROM4[2453]<=16'd57264;
ROM1[2454]<=16'd4728; ROM2[2454]<=16'd0; ROM3[2454]<=16'd23784; ROM4[2454]<=16'd57268;
ROM1[2455]<=16'd4727; ROM2[2455]<=16'd0; ROM3[2455]<=16'd23790; ROM4[2455]<=16'd57274;
ROM1[2456]<=16'd4736; ROM2[2456]<=16'd0; ROM3[2456]<=16'd23784; ROM4[2456]<=16'd57269;
ROM1[2457]<=16'd4759; ROM2[2457]<=16'd0; ROM3[2457]<=16'd23768; ROM4[2457]<=16'd57260;
ROM1[2458]<=16'd4782; ROM2[2458]<=16'd0; ROM3[2458]<=16'd23761; ROM4[2458]<=16'd57262;
ROM1[2459]<=16'd4777; ROM2[2459]<=16'd0; ROM3[2459]<=16'd23765; ROM4[2459]<=16'd57264;
ROM1[2460]<=16'd4766; ROM2[2460]<=16'd0; ROM3[2460]<=16'd23778; ROM4[2460]<=16'd57271;
ROM1[2461]<=16'd4768; ROM2[2461]<=16'd0; ROM3[2461]<=16'd23798; ROM4[2461]<=16'd57284;
ROM1[2462]<=16'd4752; ROM2[2462]<=16'd0; ROM3[2462]<=16'd23797; ROM4[2462]<=16'd57275;
ROM1[2463]<=16'd4739; ROM2[2463]<=16'd0; ROM3[2463]<=16'd23796; ROM4[2463]<=16'd57272;
ROM1[2464]<=16'd4738; ROM2[2464]<=16'd0; ROM3[2464]<=16'd23788; ROM4[2464]<=16'd57267;
ROM1[2465]<=16'd4747; ROM2[2465]<=16'd0; ROM3[2465]<=16'd23770; ROM4[2465]<=16'd57252;
ROM1[2466]<=16'd4774; ROM2[2466]<=16'd0; ROM3[2466]<=16'd23765; ROM4[2466]<=16'd57254;
ROM1[2467]<=16'd4773; ROM2[2467]<=16'd0; ROM3[2467]<=16'd23764; ROM4[2467]<=16'd57255;
ROM1[2468]<=16'd4759; ROM2[2468]<=16'd0; ROM3[2468]<=16'd23770; ROM4[2468]<=16'd57256;
ROM1[2469]<=16'd4750; ROM2[2469]<=16'd0; ROM3[2469]<=16'd23788; ROM4[2469]<=16'd57265;
ROM1[2470]<=16'd4743; ROM2[2470]<=16'd0; ROM3[2470]<=16'd23793; ROM4[2470]<=16'd57268;
ROM1[2471]<=16'd4728; ROM2[2471]<=16'd0; ROM3[2471]<=16'd23795; ROM4[2471]<=16'd57262;
ROM1[2472]<=16'd4731; ROM2[2472]<=16'd0; ROM3[2472]<=16'd23798; ROM4[2472]<=16'd57265;
ROM1[2473]<=16'd4753; ROM2[2473]<=16'd0; ROM3[2473]<=16'd23786; ROM4[2473]<=16'd57266;
ROM1[2474]<=16'd4775; ROM2[2474]<=16'd0; ROM3[2474]<=16'd23767; ROM4[2474]<=16'd57255;
ROM1[2475]<=16'd4788; ROM2[2475]<=16'd0; ROM3[2475]<=16'd23764; ROM4[2475]<=16'd57259;
ROM1[2476]<=16'd4781; ROM2[2476]<=16'd0; ROM3[2476]<=16'd23777; ROM4[2476]<=16'd57264;
ROM1[2477]<=16'd4766; ROM2[2477]<=16'd0; ROM3[2477]<=16'd23790; ROM4[2477]<=16'd57265;
ROM1[2478]<=16'd4750; ROM2[2478]<=16'd0; ROM3[2478]<=16'd23791; ROM4[2478]<=16'd57264;
ROM1[2479]<=16'd4714; ROM2[2479]<=16'd0; ROM3[2479]<=16'd23776; ROM4[2479]<=16'd57243;
ROM1[2480]<=16'd4700; ROM2[2480]<=16'd0; ROM3[2480]<=16'd23769; ROM4[2480]<=16'd57234;
ROM1[2481]<=16'd4715; ROM2[2481]<=16'd0; ROM3[2481]<=16'd23760; ROM4[2481]<=16'd57234;
ROM1[2482]<=16'd4755; ROM2[2482]<=16'd0; ROM3[2482]<=16'd23754; ROM4[2482]<=16'd57240;
ROM1[2483]<=16'd4784; ROM2[2483]<=16'd0; ROM3[2483]<=16'd23752; ROM4[2483]<=16'd57246;
ROM1[2484]<=16'd4769; ROM2[2484]<=16'd0; ROM3[2484]<=16'd23745; ROM4[2484]<=16'd57239;
ROM1[2485]<=16'd4748; ROM2[2485]<=16'd0; ROM3[2485]<=16'd23751; ROM4[2485]<=16'd57232;
ROM1[2486]<=16'd4737; ROM2[2486]<=16'd0; ROM3[2486]<=16'd23766; ROM4[2486]<=16'd57239;
ROM1[2487]<=16'd4737; ROM2[2487]<=16'd0; ROM3[2487]<=16'd23780; ROM4[2487]<=16'd57249;
ROM1[2488]<=16'd4738; ROM2[2488]<=16'd0; ROM3[2488]<=16'd23797; ROM4[2488]<=16'd57259;
ROM1[2489]<=16'd4745; ROM2[2489]<=16'd0; ROM3[2489]<=16'd23801; ROM4[2489]<=16'd57264;
ROM1[2490]<=16'd4753; ROM2[2490]<=16'd0; ROM3[2490]<=16'd23773; ROM4[2490]<=16'd57243;
ROM1[2491]<=16'd4765; ROM2[2491]<=16'd0; ROM3[2491]<=16'd23749; ROM4[2491]<=16'd57226;
ROM1[2492]<=16'd4761; ROM2[2492]<=16'd0; ROM3[2492]<=16'd23747; ROM4[2492]<=16'd57223;
ROM1[2493]<=16'd4744; ROM2[2493]<=16'd0; ROM3[2493]<=16'd23750; ROM4[2493]<=16'd57226;
ROM1[2494]<=16'd4751; ROM2[2494]<=16'd0; ROM3[2494]<=16'd23778; ROM4[2494]<=16'd57252;
ROM1[2495]<=16'd4762; ROM2[2495]<=16'd0; ROM3[2495]<=16'd23801; ROM4[2495]<=16'd57272;
ROM1[2496]<=16'd4738; ROM2[2496]<=16'd0; ROM3[2496]<=16'd23793; ROM4[2496]<=16'd57263;
ROM1[2497]<=16'd4713; ROM2[2497]<=16'd0; ROM3[2497]<=16'd23766; ROM4[2497]<=16'd57235;
ROM1[2498]<=16'd4722; ROM2[2498]<=16'd0; ROM3[2498]<=16'd23748; ROM4[2498]<=16'd57223;
ROM1[2499]<=16'd4756; ROM2[2499]<=16'd0; ROM3[2499]<=16'd23740; ROM4[2499]<=16'd57229;
ROM1[2500]<=16'd4777; ROM2[2500]<=16'd0; ROM3[2500]<=16'd23737; ROM4[2500]<=16'd57236;
ROM1[2501]<=16'd4765; ROM2[2501]<=16'd0; ROM3[2501]<=16'd23744; ROM4[2501]<=16'd57239;
ROM1[2502]<=16'd4742; ROM2[2502]<=16'd0; ROM3[2502]<=16'd23753; ROM4[2502]<=16'd57238;
ROM1[2503]<=16'd4730; ROM2[2503]<=16'd0; ROM3[2503]<=16'd23761; ROM4[2503]<=16'd57243;
ROM1[2504]<=16'd4706; ROM2[2504]<=16'd0; ROM3[2504]<=16'd23762; ROM4[2504]<=16'd57243;
ROM1[2505]<=16'd4709; ROM2[2505]<=16'd0; ROM3[2505]<=16'd23773; ROM4[2505]<=16'd57245;
ROM1[2506]<=16'd4729; ROM2[2506]<=16'd0; ROM3[2506]<=16'd23772; ROM4[2506]<=16'd57250;
ROM1[2507]<=16'd4767; ROM2[2507]<=16'd0; ROM3[2507]<=16'd23769; ROM4[2507]<=16'd57258;
ROM1[2508]<=16'd4793; ROM2[2508]<=16'd0; ROM3[2508]<=16'd23764; ROM4[2508]<=16'd57261;
ROM1[2509]<=16'd4768; ROM2[2509]<=16'd0; ROM3[2509]<=16'd23748; ROM4[2509]<=16'd57248;
ROM1[2510]<=16'd4748; ROM2[2510]<=16'd0; ROM3[2510]<=16'd23756; ROM4[2510]<=16'd57245;
ROM1[2511]<=16'd4734; ROM2[2511]<=16'd0; ROM3[2511]<=16'd23766; ROM4[2511]<=16'd57247;
ROM1[2512]<=16'd4720; ROM2[2512]<=16'd0; ROM3[2512]<=16'd23774; ROM4[2512]<=16'd57247;
ROM1[2513]<=16'd4724; ROM2[2513]<=16'd0; ROM3[2513]<=16'd23792; ROM4[2513]<=16'd57259;
ROM1[2514]<=16'd4740; ROM2[2514]<=16'd0; ROM3[2514]<=16'd23797; ROM4[2514]<=16'd57269;
ROM1[2515]<=16'd4760; ROM2[2515]<=16'd0; ROM3[2515]<=16'd23787; ROM4[2515]<=16'd57266;
ROM1[2516]<=16'd4795; ROM2[2516]<=16'd0; ROM3[2516]<=16'd23779; ROM4[2516]<=16'd57271;
ROM1[2517]<=16'd4808; ROM2[2517]<=16'd0; ROM3[2517]<=16'd23789; ROM4[2517]<=16'd57284;
ROM1[2518]<=16'd4787; ROM2[2518]<=16'd0; ROM3[2518]<=16'd23790; ROM4[2518]<=16'd57281;
ROM1[2519]<=16'd4754; ROM2[2519]<=16'd0; ROM3[2519]<=16'd23779; ROM4[2519]<=16'd57266;
ROM1[2520]<=16'd4743; ROM2[2520]<=16'd0; ROM3[2520]<=16'd23784; ROM4[2520]<=16'd57264;
ROM1[2521]<=16'd4732; ROM2[2521]<=16'd0; ROM3[2521]<=16'd23796; ROM4[2521]<=16'd57270;
ROM1[2522]<=16'd4730; ROM2[2522]<=16'd0; ROM3[2522]<=16'd23798; ROM4[2522]<=16'd57273;
ROM1[2523]<=16'd4753; ROM2[2523]<=16'd0; ROM3[2523]<=16'd23793; ROM4[2523]<=16'd57271;
ROM1[2524]<=16'd4784; ROM2[2524]<=16'd0; ROM3[2524]<=16'd23783; ROM4[2524]<=16'd57270;
ROM1[2525]<=16'd4793; ROM2[2525]<=16'd0; ROM3[2525]<=16'd23777; ROM4[2525]<=16'd57271;
ROM1[2526]<=16'd4779; ROM2[2526]<=16'd0; ROM3[2526]<=16'd23787; ROM4[2526]<=16'd57276;
ROM1[2527]<=16'd4778; ROM2[2527]<=16'd0; ROM3[2527]<=16'd23815; ROM4[2527]<=16'd57296;
ROM1[2528]<=16'd4786; ROM2[2528]<=16'd0; ROM3[2528]<=16'd23840; ROM4[2528]<=16'd57313;
ROM1[2529]<=16'd4765; ROM2[2529]<=16'd0; ROM3[2529]<=16'd23840; ROM4[2529]<=16'd57304;
ROM1[2530]<=16'd4757; ROM2[2530]<=16'd0; ROM3[2530]<=16'd23836; ROM4[2530]<=16'd57298;
ROM1[2531]<=16'd4760; ROM2[2531]<=16'd0; ROM3[2531]<=16'd23820; ROM4[2531]<=16'd57287;
ROM1[2532]<=16'd4782; ROM2[2532]<=16'd0; ROM3[2532]<=16'd23805; ROM4[2532]<=16'd57286;
ROM1[2533]<=16'd4820; ROM2[2533]<=16'd0; ROM3[2533]<=16'd23807; ROM4[2533]<=16'd57301;
ROM1[2534]<=16'd4825; ROM2[2534]<=16'd0; ROM3[2534]<=16'd23809; ROM4[2534]<=16'd57305;
ROM1[2535]<=16'd4808; ROM2[2535]<=16'd0; ROM3[2535]<=16'd23819; ROM4[2535]<=16'd57307;
ROM1[2536]<=16'd4792; ROM2[2536]<=16'd0; ROM3[2536]<=16'd23825; ROM4[2536]<=16'd57305;
ROM1[2537]<=16'd4778; ROM2[2537]<=16'd0; ROM3[2537]<=16'd23824; ROM4[2537]<=16'd57301;
ROM1[2538]<=16'd4773; ROM2[2538]<=16'd0; ROM3[2538]<=16'd23833; ROM4[2538]<=16'd57305;
ROM1[2539]<=16'd4784; ROM2[2539]<=16'd0; ROM3[2539]<=16'd23825; ROM4[2539]<=16'd57303;
ROM1[2540]<=16'd4799; ROM2[2540]<=16'd0; ROM3[2540]<=16'd23800; ROM4[2540]<=16'd57290;
ROM1[2541]<=16'd4828; ROM2[2541]<=16'd0; ROM3[2541]<=16'd23792; ROM4[2541]<=16'd57293;
ROM1[2542]<=16'd4837; ROM2[2542]<=16'd0; ROM3[2542]<=16'd23795; ROM4[2542]<=16'd57299;
ROM1[2543]<=16'd4820; ROM2[2543]<=16'd0; ROM3[2543]<=16'd23800; ROM4[2543]<=16'd57298;
ROM1[2544]<=16'd4824; ROM2[2544]<=16'd0; ROM3[2544]<=16'd23833; ROM4[2544]<=16'd57322;
ROM1[2545]<=16'd4815; ROM2[2545]<=16'd0; ROM3[2545]<=16'd23844; ROM4[2545]<=16'd57327;
ROM1[2546]<=16'd4780; ROM2[2546]<=16'd0; ROM3[2546]<=16'd23831; ROM4[2546]<=16'd57308;
ROM1[2547]<=16'd4774; ROM2[2547]<=16'd0; ROM3[2547]<=16'd23826; ROM4[2547]<=16'd57301;
ROM1[2548]<=16'd4774; ROM2[2548]<=16'd0; ROM3[2548]<=16'd23797; ROM4[2548]<=16'd57280;
ROM1[2549]<=16'd4805; ROM2[2549]<=16'd0; ROM3[2549]<=16'd23780; ROM4[2549]<=16'd57281;
ROM1[2550]<=16'd4821; ROM2[2550]<=16'd0; ROM3[2550]<=16'd23781; ROM4[2550]<=16'd57285;
ROM1[2551]<=16'd4810; ROM2[2551]<=16'd0; ROM3[2551]<=16'd23787; ROM4[2551]<=16'd57286;
ROM1[2552]<=16'd4800; ROM2[2552]<=16'd0; ROM3[2552]<=16'd23802; ROM4[2552]<=16'd57295;
ROM1[2553]<=16'd4788; ROM2[2553]<=16'd0; ROM3[2553]<=16'd23812; ROM4[2553]<=16'd57297;
ROM1[2554]<=16'd4776; ROM2[2554]<=16'd0; ROM3[2554]<=16'd23824; ROM4[2554]<=16'd57299;
ROM1[2555]<=16'd4766; ROM2[2555]<=16'd0; ROM3[2555]<=16'd23818; ROM4[2555]<=16'd57292;
ROM1[2556]<=16'd4778; ROM2[2556]<=16'd0; ROM3[2556]<=16'd23805; ROM4[2556]<=16'd57286;
ROM1[2557]<=16'd4809; ROM2[2557]<=16'd0; ROM3[2557]<=16'd23790; ROM4[2557]<=16'd57283;
ROM1[2558]<=16'd4824; ROM2[2558]<=16'd0; ROM3[2558]<=16'd23777; ROM4[2558]<=16'd57282;
ROM1[2559]<=16'd4820; ROM2[2559]<=16'd0; ROM3[2559]<=16'd23780; ROM4[2559]<=16'd57286;
ROM1[2560]<=16'd4814; ROM2[2560]<=16'd0; ROM3[2560]<=16'd23795; ROM4[2560]<=16'd57294;
ROM1[2561]<=16'd4812; ROM2[2561]<=16'd0; ROM3[2561]<=16'd23819; ROM4[2561]<=16'd57306;
ROM1[2562]<=16'd4785; ROM2[2562]<=16'd0; ROM3[2562]<=16'd23817; ROM4[2562]<=16'd57300;
ROM1[2563]<=16'd4764; ROM2[2563]<=16'd0; ROM3[2563]<=16'd23812; ROM4[2563]<=16'd57290;
ROM1[2564]<=16'd4763; ROM2[2564]<=16'd0; ROM3[2564]<=16'd23810; ROM4[2564]<=16'd57283;
ROM1[2565]<=16'd4775; ROM2[2565]<=16'd0; ROM3[2565]<=16'd23790; ROM4[2565]<=16'd57276;
ROM1[2566]<=16'd4809; ROM2[2566]<=16'd0; ROM3[2566]<=16'd23779; ROM4[2566]<=16'd57282;
ROM1[2567]<=16'd4818; ROM2[2567]<=16'd0; ROM3[2567]<=16'd23789; ROM4[2567]<=16'd57292;
ROM1[2568]<=16'd4804; ROM2[2568]<=16'd0; ROM3[2568]<=16'd23798; ROM4[2568]<=16'd57293;
ROM1[2569]<=16'd4792; ROM2[2569]<=16'd0; ROM3[2569]<=16'd23808; ROM4[2569]<=16'd57294;
ROM1[2570]<=16'd4785; ROM2[2570]<=16'd0; ROM3[2570]<=16'd23822; ROM4[2570]<=16'd57299;
ROM1[2571]<=16'd4770; ROM2[2571]<=16'd0; ROM3[2571]<=16'd23834; ROM4[2571]<=16'd57299;
ROM1[2572]<=16'd4758; ROM2[2572]<=16'd0; ROM3[2572]<=16'd23825; ROM4[2572]<=16'd57288;
ROM1[2573]<=16'd4770; ROM2[2573]<=16'd0; ROM3[2573]<=16'd23809; ROM4[2573]<=16'd57285;
ROM1[2574]<=16'd4810; ROM2[2574]<=16'd0; ROM3[2574]<=16'd23805; ROM4[2574]<=16'd57288;
ROM1[2575]<=16'd4827; ROM2[2575]<=16'd0; ROM3[2575]<=16'd23804; ROM4[2575]<=16'd57294;
ROM1[2576]<=16'd4821; ROM2[2576]<=16'd0; ROM3[2576]<=16'd23812; ROM4[2576]<=16'd57302;
ROM1[2577]<=16'd4800; ROM2[2577]<=16'd0; ROM3[2577]<=16'd23817; ROM4[2577]<=16'd57297;
ROM1[2578]<=16'd4783; ROM2[2578]<=16'd0; ROM3[2578]<=16'd23817; ROM4[2578]<=16'd57295;
ROM1[2579]<=16'd4761; ROM2[2579]<=16'd0; ROM3[2579]<=16'd23814; ROM4[2579]<=16'd57291;
ROM1[2580]<=16'd4749; ROM2[2580]<=16'd0; ROM3[2580]<=16'd23808; ROM4[2580]<=16'd57285;
ROM1[2581]<=16'd4769; ROM2[2581]<=16'd0; ROM3[2581]<=16'd23806; ROM4[2581]<=16'd57289;
ROM1[2582]<=16'd4814; ROM2[2582]<=16'd0; ROM3[2582]<=16'd23805; ROM4[2582]<=16'd57297;
ROM1[2583]<=16'd4844; ROM2[2583]<=16'd0; ROM3[2583]<=16'd23800; ROM4[2583]<=16'd57305;
ROM1[2584]<=16'd4837; ROM2[2584]<=16'd0; ROM3[2584]<=16'd23807; ROM4[2584]<=16'd57310;
ROM1[2585]<=16'd4822; ROM2[2585]<=16'd0; ROM3[2585]<=16'd23819; ROM4[2585]<=16'd57315;
ROM1[2586]<=16'd4810; ROM2[2586]<=16'd0; ROM3[2586]<=16'd23832; ROM4[2586]<=16'd57324;
ROM1[2587]<=16'd4797; ROM2[2587]<=16'd0; ROM3[2587]<=16'd23841; ROM4[2587]<=16'd57322;
ROM1[2588]<=16'd4783; ROM2[2588]<=16'd0; ROM3[2588]<=16'd23844; ROM4[2588]<=16'd57321;
ROM1[2589]<=16'd4780; ROM2[2589]<=16'd0; ROM3[2589]<=16'd23835; ROM4[2589]<=16'd57315;
ROM1[2590]<=16'd4797; ROM2[2590]<=16'd0; ROM3[2590]<=16'd23813; ROM4[2590]<=16'd57302;
ROM1[2591]<=16'd4823; ROM2[2591]<=16'd0; ROM3[2591]<=16'd23798; ROM4[2591]<=16'd57298;
ROM1[2592]<=16'd4821; ROM2[2592]<=16'd0; ROM3[2592]<=16'd23790; ROM4[2592]<=16'd57294;
ROM1[2593]<=16'd4803; ROM2[2593]<=16'd0; ROM3[2593]<=16'd23793; ROM4[2593]<=16'd57292;
ROM1[2594]<=16'd4783; ROM2[2594]<=16'd0; ROM3[2594]<=16'd23796; ROM4[2594]<=16'd57292;
ROM1[2595]<=16'd4781; ROM2[2595]<=16'd0; ROM3[2595]<=16'd23811; ROM4[2595]<=16'd57303;
ROM1[2596]<=16'd4776; ROM2[2596]<=16'd0; ROM3[2596]<=16'd23818; ROM4[2596]<=16'd57308;
ROM1[2597]<=16'd4769; ROM2[2597]<=16'd0; ROM3[2597]<=16'd23804; ROM4[2597]<=16'd57294;
ROM1[2598]<=16'd4785; ROM2[2598]<=16'd0; ROM3[2598]<=16'd23793; ROM4[2598]<=16'd57287;
ROM1[2599]<=16'd4803; ROM2[2599]<=16'd0; ROM3[2599]<=16'd23768; ROM4[2599]<=16'd57274;
ROM1[2600]<=16'd4801; ROM2[2600]<=16'd0; ROM3[2600]<=16'd23758; ROM4[2600]<=16'd57267;
ROM1[2601]<=16'd4795; ROM2[2601]<=16'd0; ROM3[2601]<=16'd23774; ROM4[2601]<=16'd57273;
ROM1[2602]<=16'd4782; ROM2[2602]<=16'd0; ROM3[2602]<=16'd23793; ROM4[2602]<=16'd57278;
ROM1[2603]<=16'd4765; ROM2[2603]<=16'd0; ROM3[2603]<=16'd23794; ROM4[2603]<=16'd57274;
ROM1[2604]<=16'd4759; ROM2[2604]<=16'd0; ROM3[2604]<=16'd23805; ROM4[2604]<=16'd57281;
ROM1[2605]<=16'd4765; ROM2[2605]<=16'd0; ROM3[2605]<=16'd23822; ROM4[2605]<=16'd57292;
ROM1[2606]<=16'd4775; ROM2[2606]<=16'd0; ROM3[2606]<=16'd23818; ROM4[2606]<=16'd57294;
ROM1[2607]<=16'd4799; ROM2[2607]<=16'd0; ROM3[2607]<=16'd23805; ROM4[2607]<=16'd57294;
ROM1[2608]<=16'd4823; ROM2[2608]<=16'd0; ROM3[2608]<=16'd23800; ROM4[2608]<=16'd57297;
ROM1[2609]<=16'd4825; ROM2[2609]<=16'd0; ROM3[2609]<=16'd23814; ROM4[2609]<=16'd57313;
ROM1[2610]<=16'd4806; ROM2[2610]<=16'd0; ROM3[2610]<=16'd23821; ROM4[2610]<=16'd57314;
ROM1[2611]<=16'd4771; ROM2[2611]<=16'd0; ROM3[2611]<=16'd23811; ROM4[2611]<=16'd57296;
ROM1[2612]<=16'd4749; ROM2[2612]<=16'd0; ROM3[2612]<=16'd23814; ROM4[2612]<=16'd57293;
ROM1[2613]<=16'd4732; ROM2[2613]<=16'd0; ROM3[2613]<=16'd23805; ROM4[2613]<=16'd57281;
ROM1[2614]<=16'd4744; ROM2[2614]<=16'd0; ROM3[2614]<=16'd23803; ROM4[2614]<=16'd57278;
ROM1[2615]<=16'd4789; ROM2[2615]<=16'd0; ROM3[2615]<=16'd23818; ROM4[2615]<=16'd57297;
ROM1[2616]<=16'd4803; ROM2[2616]<=16'd0; ROM3[2616]<=16'd23792; ROM4[2616]<=16'd57281;
ROM1[2617]<=16'd4792; ROM2[2617]<=16'd0; ROM3[2617]<=16'd23772; ROM4[2617]<=16'd57263;
ROM1[2618]<=16'd4780; ROM2[2618]<=16'd0; ROM3[2618]<=16'd23774; ROM4[2618]<=16'd57260;
ROM1[2619]<=16'd4766; ROM2[2619]<=16'd0; ROM3[2619]<=16'd23779; ROM4[2619]<=16'd57258;
ROM1[2620]<=16'd4765; ROM2[2620]<=16'd0; ROM3[2620]<=16'd23793; ROM4[2620]<=16'd57268;
ROM1[2621]<=16'd4748; ROM2[2621]<=16'd0; ROM3[2621]<=16'd23800; ROM4[2621]<=16'd57268;
ROM1[2622]<=16'd4744; ROM2[2622]<=16'd0; ROM3[2622]<=16'd23801; ROM4[2622]<=16'd57271;
ROM1[2623]<=16'd4771; ROM2[2623]<=16'd0; ROM3[2623]<=16'd23795; ROM4[2623]<=16'd57276;
ROM1[2624]<=16'd4807; ROM2[2624]<=16'd0; ROM3[2624]<=16'd23784; ROM4[2624]<=16'd57274;
ROM1[2625]<=16'd4818; ROM2[2625]<=16'd0; ROM3[2625]<=16'd23779; ROM4[2625]<=16'd57274;
ROM1[2626]<=16'd4800; ROM2[2626]<=16'd0; ROM3[2626]<=16'd23782; ROM4[2626]<=16'd57270;
ROM1[2627]<=16'd4783; ROM2[2627]<=16'd0; ROM3[2627]<=16'd23793; ROM4[2627]<=16'd57270;
ROM1[2628]<=16'd4783; ROM2[2628]<=16'd0; ROM3[2628]<=16'd23810; ROM4[2628]<=16'd57286;
ROM1[2629]<=16'd4766; ROM2[2629]<=16'd0; ROM3[2629]<=16'd23815; ROM4[2629]<=16'd57283;
ROM1[2630]<=16'd4749; ROM2[2630]<=16'd0; ROM3[2630]<=16'd23797; ROM4[2630]<=16'd57267;
ROM1[2631]<=16'd4761; ROM2[2631]<=16'd0; ROM3[2631]<=16'd23787; ROM4[2631]<=16'd57265;
ROM1[2632]<=16'd4788; ROM2[2632]<=16'd0; ROM3[2632]<=16'd23774; ROM4[2632]<=16'd57261;
ROM1[2633]<=16'd4804; ROM2[2633]<=16'd0; ROM3[2633]<=16'd23764; ROM4[2633]<=16'd57260;
ROM1[2634]<=16'd4791; ROM2[2634]<=16'd0; ROM3[2634]<=16'd23765; ROM4[2634]<=16'd57259;
ROM1[2635]<=16'd4758; ROM2[2635]<=16'd0; ROM3[2635]<=16'd23762; ROM4[2635]<=16'd57246;
ROM1[2636]<=16'd4746; ROM2[2636]<=16'd0; ROM3[2636]<=16'd23773; ROM4[2636]<=16'd57252;
ROM1[2637]<=16'd4745; ROM2[2637]<=16'd0; ROM3[2637]<=16'd23791; ROM4[2637]<=16'd57267;
ROM1[2638]<=16'd4739; ROM2[2638]<=16'd0; ROM3[2638]<=16'd23799; ROM4[2638]<=16'd57272;
ROM1[2639]<=16'd4747; ROM2[2639]<=16'd0; ROM3[2639]<=16'd23802; ROM4[2639]<=16'd57279;
ROM1[2640]<=16'd4766; ROM2[2640]<=16'd0; ROM3[2640]<=16'd23788; ROM4[2640]<=16'd57269;
ROM1[2641]<=16'd4792; ROM2[2641]<=16'd0; ROM3[2641]<=16'd23769; ROM4[2641]<=16'd57263;
ROM1[2642]<=16'd4802; ROM2[2642]<=16'd0; ROM3[2642]<=16'd23769; ROM4[2642]<=16'd57270;
ROM1[2643]<=16'd4790; ROM2[2643]<=16'd0; ROM3[2643]<=16'd23777; ROM4[2643]<=16'd57275;
ROM1[2644]<=16'd4776; ROM2[2644]<=16'd0; ROM3[2644]<=16'd23786; ROM4[2644]<=16'd57278;
ROM1[2645]<=16'd4770; ROM2[2645]<=16'd0; ROM3[2645]<=16'd23796; ROM4[2645]<=16'd57285;
ROM1[2646]<=16'd4758; ROM2[2646]<=16'd0; ROM3[2646]<=16'd23799; ROM4[2646]<=16'd57286;
ROM1[2647]<=16'd4757; ROM2[2647]<=16'd0; ROM3[2647]<=16'd23794; ROM4[2647]<=16'd57281;
ROM1[2648]<=16'd4778; ROM2[2648]<=16'd0; ROM3[2648]<=16'd23788; ROM4[2648]<=16'd57281;
ROM1[2649]<=16'd4800; ROM2[2649]<=16'd0; ROM3[2649]<=16'd23767; ROM4[2649]<=16'd57273;
ROM1[2650]<=16'd4797; ROM2[2650]<=16'd0; ROM3[2650]<=16'd23756; ROM4[2650]<=16'd57266;
ROM1[2651]<=16'd4786; ROM2[2651]<=16'd0; ROM3[2651]<=16'd23766; ROM4[2651]<=16'd57275;
ROM1[2652]<=16'd4770; ROM2[2652]<=16'd0; ROM3[2652]<=16'd23773; ROM4[2652]<=16'd57277;
ROM1[2653]<=16'd4755; ROM2[2653]<=16'd0; ROM3[2653]<=16'd23782; ROM4[2653]<=16'd57279;
ROM1[2654]<=16'd4742; ROM2[2654]<=16'd0; ROM3[2654]<=16'd23793; ROM4[2654]<=16'd57287;
ROM1[2655]<=16'd4744; ROM2[2655]<=16'd0; ROM3[2655]<=16'd23805; ROM4[2655]<=16'd57289;
ROM1[2656]<=16'd4765; ROM2[2656]<=16'd0; ROM3[2656]<=16'd23802; ROM4[2656]<=16'd57292;
ROM1[2657]<=16'd4788; ROM2[2657]<=16'd0; ROM3[2657]<=16'd23784; ROM4[2657]<=16'd57285;
ROM1[2658]<=16'd4818; ROM2[2658]<=16'd0; ROM3[2658]<=16'd23785; ROM4[2658]<=16'd57294;
ROM1[2659]<=16'd4812; ROM2[2659]<=16'd0; ROM3[2659]<=16'd23786; ROM4[2659]<=16'd57294;
ROM1[2660]<=16'd4772; ROM2[2660]<=16'd0; ROM3[2660]<=16'd23772; ROM4[2660]<=16'd57273;
ROM1[2661]<=16'd4757; ROM2[2661]<=16'd0; ROM3[2661]<=16'd23782; ROM4[2661]<=16'd57273;
ROM1[2662]<=16'd4747; ROM2[2662]<=16'd0; ROM3[2662]<=16'd23788; ROM4[2662]<=16'd57273;
ROM1[2663]<=16'd4734; ROM2[2663]<=16'd0; ROM3[2663]<=16'd23787; ROM4[2663]<=16'd57267;
ROM1[2664]<=16'd4748; ROM2[2664]<=16'd0; ROM3[2664]<=16'd23794; ROM4[2664]<=16'd57276;
ROM1[2665]<=16'd4786; ROM2[2665]<=16'd0; ROM3[2665]<=16'd23792; ROM4[2665]<=16'd57282;
ROM1[2666]<=16'd4816; ROM2[2666]<=16'd0; ROM3[2666]<=16'd23782; ROM4[2666]<=16'd57283;
ROM1[2667]<=16'd4818; ROM2[2667]<=16'd0; ROM3[2667]<=16'd23786; ROM4[2667]<=16'd57290;
ROM1[2668]<=16'd4807; ROM2[2668]<=16'd0; ROM3[2668]<=16'd23801; ROM4[2668]<=16'd57299;
ROM1[2669]<=16'd4782; ROM2[2669]<=16'd0; ROM3[2669]<=16'd23807; ROM4[2669]<=16'd57290;
ROM1[2670]<=16'd4768; ROM2[2670]<=16'd0; ROM3[2670]<=16'd23812; ROM4[2670]<=16'd57287;
ROM1[2671]<=16'd4760; ROM2[2671]<=16'd0; ROM3[2671]<=16'd23815; ROM4[2671]<=16'd57285;
ROM1[2672]<=16'd4762; ROM2[2672]<=16'd0; ROM3[2672]<=16'd23809; ROM4[2672]<=16'd57281;
ROM1[2673]<=16'd4788; ROM2[2673]<=16'd0; ROM3[2673]<=16'd23800; ROM4[2673]<=16'd57284;
ROM1[2674]<=16'd4814; ROM2[2674]<=16'd0; ROM3[2674]<=16'd23780; ROM4[2674]<=16'd57279;
ROM1[2675]<=16'd4812; ROM2[2675]<=16'd0; ROM3[2675]<=16'd23765; ROM4[2675]<=16'd57273;
ROM1[2676]<=16'd4800; ROM2[2676]<=16'd0; ROM3[2676]<=16'd23770; ROM4[2676]<=16'd57274;
ROM1[2677]<=16'd4789; ROM2[2677]<=16'd0; ROM3[2677]<=16'd23782; ROM4[2677]<=16'd57277;
ROM1[2678]<=16'd4777; ROM2[2678]<=16'd0; ROM3[2678]<=16'd23786; ROM4[2678]<=16'd57276;
ROM1[2679]<=16'd4759; ROM2[2679]<=16'd0; ROM3[2679]<=16'd23785; ROM4[2679]<=16'd57266;
ROM1[2680]<=16'd4752; ROM2[2680]<=16'd0; ROM3[2680]<=16'd23776; ROM4[2680]<=16'd57261;
ROM1[2681]<=16'd4761; ROM2[2681]<=16'd0; ROM3[2681]<=16'd23762; ROM4[2681]<=16'd57254;
ROM1[2682]<=16'd4783; ROM2[2682]<=16'd0; ROM3[2682]<=16'd23734; ROM4[2682]<=16'd57242;
ROM1[2683]<=16'd4800; ROM2[2683]<=16'd0; ROM3[2683]<=16'd23721; ROM4[2683]<=16'd57242;
ROM1[2684]<=16'd4792; ROM2[2684]<=16'd0; ROM3[2684]<=16'd23724; ROM4[2684]<=16'd57243;
ROM1[2685]<=16'd4769; ROM2[2685]<=16'd0; ROM3[2685]<=16'd23720; ROM4[2685]<=16'd57234;
ROM1[2686]<=16'd4761; ROM2[2686]<=16'd0; ROM3[2686]<=16'd23736; ROM4[2686]<=16'd57241;
ROM1[2687]<=16'd4760; ROM2[2687]<=16'd0; ROM3[2687]<=16'd23752; ROM4[2687]<=16'd57256;
ROM1[2688]<=16'd4751; ROM2[2688]<=16'd0; ROM3[2688]<=16'd23752; ROM4[2688]<=16'd57258;
ROM1[2689]<=16'd4757; ROM2[2689]<=16'd0; ROM3[2689]<=16'd23749; ROM4[2689]<=16'd57257;
ROM1[2690]<=16'd4781; ROM2[2690]<=16'd0; ROM3[2690]<=16'd23737; ROM4[2690]<=16'd57254;
ROM1[2691]<=16'd4801; ROM2[2691]<=16'd0; ROM3[2691]<=16'd23723; ROM4[2691]<=16'd57248;
ROM1[2692]<=16'd4789; ROM2[2692]<=16'd0; ROM3[2692]<=16'd23718; ROM4[2692]<=16'd57240;
ROM1[2693]<=16'd4782; ROM2[2693]<=16'd0; ROM3[2693]<=16'd23740; ROM4[2693]<=16'd57253;
ROM1[2694]<=16'd4774; ROM2[2694]<=16'd0; ROM3[2694]<=16'd23762; ROM4[2694]<=16'd57266;
ROM1[2695]<=16'd4748; ROM2[2695]<=16'd0; ROM3[2695]<=16'd23757; ROM4[2695]<=16'd57254;
ROM1[2696]<=16'd4736; ROM2[2696]<=16'd0; ROM3[2696]<=16'd23762; ROM4[2696]<=16'd57255;
ROM1[2697]<=16'd4736; ROM2[2697]<=16'd0; ROM3[2697]<=16'd23761; ROM4[2697]<=16'd57254;
ROM1[2698]<=16'd4745; ROM2[2698]<=16'd0; ROM3[2698]<=16'd23742; ROM4[2698]<=16'd57241;
ROM1[2699]<=16'd4788; ROM2[2699]<=16'd0; ROM3[2699]<=16'd23738; ROM4[2699]<=16'd57252;
ROM1[2700]<=16'd4824; ROM2[2700]<=16'd0; ROM3[2700]<=16'd23755; ROM4[2700]<=16'd57279;
ROM1[2701]<=16'd4816; ROM2[2701]<=16'd0; ROM3[2701]<=16'd23761; ROM4[2701]<=16'd57281;
ROM1[2702]<=16'd4776; ROM2[2702]<=16'd0; ROM3[2702]<=16'd23748; ROM4[2702]<=16'd57262;
ROM1[2703]<=16'd4748; ROM2[2703]<=16'd0; ROM3[2703]<=16'd23747; ROM4[2703]<=16'd57252;
ROM1[2704]<=16'd4721; ROM2[2704]<=16'd0; ROM3[2704]<=16'd23750; ROM4[2704]<=16'd57247;
ROM1[2705]<=16'd4711; ROM2[2705]<=16'd0; ROM3[2705]<=16'd23750; ROM4[2705]<=16'd57245;
ROM1[2706]<=16'd4739; ROM2[2706]<=16'd0; ROM3[2706]<=16'd23756; ROM4[2706]<=16'd57258;
ROM1[2707]<=16'd4793; ROM2[2707]<=16'd0; ROM3[2707]<=16'd23765; ROM4[2707]<=16'd57281;
ROM1[2708]<=16'd4806; ROM2[2708]<=16'd0; ROM3[2708]<=16'd23752; ROM4[2708]<=16'd57276;
ROM1[2709]<=16'd4770; ROM2[2709]<=16'd0; ROM3[2709]<=16'd23735; ROM4[2709]<=16'd57250;
ROM1[2710]<=16'd4753; ROM2[2710]<=16'd0; ROM3[2710]<=16'd23749; ROM4[2710]<=16'd57256;
ROM1[2711]<=16'd4734; ROM2[2711]<=16'd0; ROM3[2711]<=16'd23755; ROM4[2711]<=16'd57252;
ROM1[2712]<=16'd4708; ROM2[2712]<=16'd0; ROM3[2712]<=16'd23751; ROM4[2712]<=16'd57242;
ROM1[2713]<=16'd4711; ROM2[2713]<=16'd0; ROM3[2713]<=16'd23768; ROM4[2713]<=16'd57255;
ROM1[2714]<=16'd4740; ROM2[2714]<=16'd0; ROM3[2714]<=16'd23784; ROM4[2714]<=16'd57273;
ROM1[2715]<=16'd4769; ROM2[2715]<=16'd0; ROM3[2715]<=16'd23773; ROM4[2715]<=16'd57276;
ROM1[2716]<=16'd4787; ROM2[2716]<=16'd0; ROM3[2716]<=16'd23750; ROM4[2716]<=16'd57262;
ROM1[2717]<=16'd4795; ROM2[2717]<=16'd0; ROM3[2717]<=16'd23751; ROM4[2717]<=16'd57272;
ROM1[2718]<=16'd4779; ROM2[2718]<=16'd0; ROM3[2718]<=16'd23754; ROM4[2718]<=16'd57271;
ROM1[2719]<=16'd4763; ROM2[2719]<=16'd0; ROM3[2719]<=16'd23757; ROM4[2719]<=16'd57266;
ROM1[2720]<=16'd4750; ROM2[2720]<=16'd0; ROM3[2720]<=16'd23766; ROM4[2720]<=16'd57269;
ROM1[2721]<=16'd4728; ROM2[2721]<=16'd0; ROM3[2721]<=16'd23769; ROM4[2721]<=16'd57267;
ROM1[2722]<=16'd4725; ROM2[2722]<=16'd0; ROM3[2722]<=16'd23762; ROM4[2722]<=16'd57260;
ROM1[2723]<=16'd4744; ROM2[2723]<=16'd0; ROM3[2723]<=16'd23752; ROM4[2723]<=16'd57257;
ROM1[2724]<=16'd4784; ROM2[2724]<=16'd0; ROM3[2724]<=16'd23747; ROM4[2724]<=16'd57264;
ROM1[2725]<=16'd4795; ROM2[2725]<=16'd0; ROM3[2725]<=16'd23745; ROM4[2725]<=16'd57267;
ROM1[2726]<=16'd4783; ROM2[2726]<=16'd0; ROM3[2726]<=16'd23758; ROM4[2726]<=16'd57274;
ROM1[2727]<=16'd4765; ROM2[2727]<=16'd0; ROM3[2727]<=16'd23777; ROM4[2727]<=16'd57280;
ROM1[2728]<=16'd4758; ROM2[2728]<=16'd0; ROM3[2728]<=16'd23789; ROM4[2728]<=16'd57287;
ROM1[2729]<=16'd4750; ROM2[2729]<=16'd0; ROM3[2729]<=16'd23795; ROM4[2729]<=16'd57284;
ROM1[2730]<=16'd4732; ROM2[2730]<=16'd0; ROM3[2730]<=16'd23782; ROM4[2730]<=16'd57267;
ROM1[2731]<=16'd4742; ROM2[2731]<=16'd0; ROM3[2731]<=16'd23766; ROM4[2731]<=16'd57261;
ROM1[2732]<=16'd4784; ROM2[2732]<=16'd0; ROM3[2732]<=16'd23759; ROM4[2732]<=16'd57266;
ROM1[2733]<=16'd4809; ROM2[2733]<=16'd0; ROM3[2733]<=16'd23755; ROM4[2733]<=16'd57272;
ROM1[2734]<=16'd4801; ROM2[2734]<=16'd0; ROM3[2734]<=16'd23759; ROM4[2734]<=16'd57277;
ROM1[2735]<=16'd4793; ROM2[2735]<=16'd0; ROM3[2735]<=16'd23773; ROM4[2735]<=16'd57283;
ROM1[2736]<=16'd4776; ROM2[2736]<=16'd0; ROM3[2736]<=16'd23783; ROM4[2736]<=16'd57281;
ROM1[2737]<=16'd4758; ROM2[2737]<=16'd0; ROM3[2737]<=16'd23786; ROM4[2737]<=16'd57277;
ROM1[2738]<=16'd4751; ROM2[2738]<=16'd0; ROM3[2738]<=16'd23790; ROM4[2738]<=16'd57279;
ROM1[2739]<=16'd4752; ROM2[2739]<=16'd0; ROM3[2739]<=16'd23786; ROM4[2739]<=16'd57277;
ROM1[2740]<=16'd4776; ROM2[2740]<=16'd0; ROM3[2740]<=16'd23777; ROM4[2740]<=16'd57278;
ROM1[2741]<=16'd4810; ROM2[2741]<=16'd0; ROM3[2741]<=16'd23771; ROM4[2741]<=16'd57285;
ROM1[2742]<=16'd4812; ROM2[2742]<=16'd0; ROM3[2742]<=16'd23771; ROM4[2742]<=16'd57285;
ROM1[2743]<=16'd4791; ROM2[2743]<=16'd0; ROM3[2743]<=16'd23771; ROM4[2743]<=16'd57284;
ROM1[2744]<=16'd4779; ROM2[2744]<=16'd0; ROM3[2744]<=16'd23781; ROM4[2744]<=16'd57290;
ROM1[2745]<=16'd4769; ROM2[2745]<=16'd0; ROM3[2745]<=16'd23794; ROM4[2745]<=16'd57298;
ROM1[2746]<=16'd4764; ROM2[2746]<=16'd0; ROM3[2746]<=16'd23809; ROM4[2746]<=16'd57311;
ROM1[2747]<=16'd4778; ROM2[2747]<=16'd0; ROM3[2747]<=16'd23821; ROM4[2747]<=16'd57319;
ROM1[2748]<=16'd4789; ROM2[2748]<=16'd0; ROM3[2748]<=16'd23810; ROM4[2748]<=16'd57312;
ROM1[2749]<=16'd4814; ROM2[2749]<=16'd0; ROM3[2749]<=16'd23794; ROM4[2749]<=16'd57310;
ROM1[2750]<=16'd4825; ROM2[2750]<=16'd0; ROM3[2750]<=16'd23800; ROM4[2750]<=16'd57321;
ROM1[2751]<=16'd4817; ROM2[2751]<=16'd0; ROM3[2751]<=16'd23816; ROM4[2751]<=16'd57337;
ROM1[2752]<=16'd4805; ROM2[2752]<=16'd0; ROM3[2752]<=16'd23819; ROM4[2752]<=16'd57340;
ROM1[2753]<=16'd4789; ROM2[2753]<=16'd0; ROM3[2753]<=16'd23810; ROM4[2753]<=16'd57328;
ROM1[2754]<=16'd4779; ROM2[2754]<=16'd0; ROM3[2754]<=16'd23815; ROM4[2754]<=16'd57326;
ROM1[2755]<=16'd4763; ROM2[2755]<=16'd0; ROM3[2755]<=16'd23805; ROM4[2755]<=16'd57315;
ROM1[2756]<=16'd4760; ROM2[2756]<=16'd0; ROM3[2756]<=16'd23783; ROM4[2756]<=16'd57300;
ROM1[2757]<=16'd4789; ROM2[2757]<=16'd0; ROM3[2757]<=16'd23771; ROM4[2757]<=16'd57301;
ROM1[2758]<=16'd4814; ROM2[2758]<=16'd0; ROM3[2758]<=16'd23763; ROM4[2758]<=16'd57302;
ROM1[2759]<=16'd4827; ROM2[2759]<=16'd0; ROM3[2759]<=16'd23781; ROM4[2759]<=16'd57315;
ROM1[2760]<=16'd4807; ROM2[2760]<=16'd0; ROM3[2760]<=16'd23790; ROM4[2760]<=16'd57316;
ROM1[2761]<=16'd4769; ROM2[2761]<=16'd0; ROM3[2761]<=16'd23780; ROM4[2761]<=16'd57298;
ROM1[2762]<=16'd4741; ROM2[2762]<=16'd0; ROM3[2762]<=16'd23770; ROM4[2762]<=16'd57286;
ROM1[2763]<=16'd4722; ROM2[2763]<=16'd0; ROM3[2763]<=16'd23762; ROM4[2763]<=16'd57274;
ROM1[2764]<=16'd4731; ROM2[2764]<=16'd0; ROM3[2764]<=16'd23758; ROM4[2764]<=16'd57272;
ROM1[2765]<=16'd4767; ROM2[2765]<=16'd0; ROM3[2765]<=16'd23756; ROM4[2765]<=16'd57279;
ROM1[2766]<=16'd4790; ROM2[2766]<=16'd0; ROM3[2766]<=16'd23740; ROM4[2766]<=16'd57272;
ROM1[2767]<=16'd4773; ROM2[2767]<=16'd0; ROM3[2767]<=16'd23724; ROM4[2767]<=16'd57255;
ROM1[2768]<=16'd4764; ROM2[2768]<=16'd0; ROM3[2768]<=16'd23735; ROM4[2768]<=16'd57264;
ROM1[2769]<=16'd4757; ROM2[2769]<=16'd0; ROM3[2769]<=16'd23754; ROM4[2769]<=16'd57275;
ROM1[2770]<=16'd4734; ROM2[2770]<=16'd0; ROM3[2770]<=16'd23760; ROM4[2770]<=16'd57269;
ROM1[2771]<=16'd4713; ROM2[2771]<=16'd0; ROM3[2771]<=16'd23761; ROM4[2771]<=16'd57262;
ROM1[2772]<=16'd4713; ROM2[2772]<=16'd0; ROM3[2772]<=16'd23762; ROM4[2772]<=16'd57259;
ROM1[2773]<=16'd4736; ROM2[2773]<=16'd0; ROM3[2773]<=16'd23752; ROM4[2773]<=16'd57259;
ROM1[2774]<=16'd4764; ROM2[2774]<=16'd0; ROM3[2774]<=16'd23738; ROM4[2774]<=16'd57255;
ROM1[2775]<=16'd4772; ROM2[2775]<=16'd0; ROM3[2775]<=16'd23736; ROM4[2775]<=16'd57255;
ROM1[2776]<=16'd4772; ROM2[2776]<=16'd0; ROM3[2776]<=16'd23750; ROM4[2776]<=16'd57264;
ROM1[2777]<=16'd4760; ROM2[2777]<=16'd0; ROM3[2777]<=16'd23765; ROM4[2777]<=16'd57267;
ROM1[2778]<=16'd4748; ROM2[2778]<=16'd0; ROM3[2778]<=16'd23769; ROM4[2778]<=16'd57266;
ROM1[2779]<=16'd4737; ROM2[2779]<=16'd0; ROM3[2779]<=16'd23777; ROM4[2779]<=16'd57268;
ROM1[2780]<=16'd4728; ROM2[2780]<=16'd0; ROM3[2780]<=16'd23777; ROM4[2780]<=16'd57265;
ROM1[2781]<=16'd4737; ROM2[2781]<=16'd0; ROM3[2781]<=16'd23773; ROM4[2781]<=16'd57265;
ROM1[2782]<=16'd4774; ROM2[2782]<=16'd0; ROM3[2782]<=16'd23767; ROM4[2782]<=16'd57271;
ROM1[2783]<=16'd4808; ROM2[2783]<=16'd0; ROM3[2783]<=16'd23768; ROM4[2783]<=16'd57284;
ROM1[2784]<=16'd4820; ROM2[2784]<=16'd0; ROM3[2784]<=16'd23786; ROM4[2784]<=16'd57297;
ROM1[2785]<=16'd4795; ROM2[2785]<=16'd0; ROM3[2785]<=16'd23782; ROM4[2785]<=16'd57285;
ROM1[2786]<=16'd4773; ROM2[2786]<=16'd0; ROM3[2786]<=16'd23780; ROM4[2786]<=16'd57274;
ROM1[2787]<=16'd4769; ROM2[2787]<=16'd0; ROM3[2787]<=16'd23794; ROM4[2787]<=16'd57284;
ROM1[2788]<=16'd4755; ROM2[2788]<=16'd0; ROM3[2788]<=16'd23792; ROM4[2788]<=16'd57281;
ROM1[2789]<=16'd4773; ROM2[2789]<=16'd0; ROM3[2789]<=16'd23800; ROM4[2789]<=16'd57293;
ROM1[2790]<=16'd4831; ROM2[2790]<=16'd0; ROM3[2790]<=16'd23824; ROM4[2790]<=16'd57326;
ROM1[2791]<=16'd4856; ROM2[2791]<=16'd0; ROM3[2791]<=16'd23809; ROM4[2791]<=16'd57324;
ROM1[2792]<=16'd4833; ROM2[2792]<=16'd0; ROM3[2792]<=16'd23780; ROM4[2792]<=16'd57300;
ROM1[2793]<=16'd4808; ROM2[2793]<=16'd0; ROM3[2793]<=16'd23781; ROM4[2793]<=16'd57294;
ROM1[2794]<=16'd4783; ROM2[2794]<=16'd0; ROM3[2794]<=16'd23780; ROM4[2794]<=16'd57287;
ROM1[2795]<=16'd4770; ROM2[2795]<=16'd0; ROM3[2795]<=16'd23785; ROM4[2795]<=16'd57289;
ROM1[2796]<=16'd4766; ROM2[2796]<=16'd0; ROM3[2796]<=16'd23802; ROM4[2796]<=16'd57300;
ROM1[2797]<=16'd4774; ROM2[2797]<=16'd0; ROM3[2797]<=16'd23803; ROM4[2797]<=16'd57301;
ROM1[2798]<=16'd4792; ROM2[2798]<=16'd0; ROM3[2798]<=16'd23785; ROM4[2798]<=16'd57292;
ROM1[2799]<=16'd4815; ROM2[2799]<=16'd0; ROM3[2799]<=16'd23767; ROM4[2799]<=16'd57283;
ROM1[2800]<=16'd4821; ROM2[2800]<=16'd0; ROM3[2800]<=16'd23771; ROM4[2800]<=16'd57291;
ROM1[2801]<=16'd4815; ROM2[2801]<=16'd0; ROM3[2801]<=16'd23792; ROM4[2801]<=16'd57305;
ROM1[2802]<=16'd4803; ROM2[2802]<=16'd0; ROM3[2802]<=16'd23806; ROM4[2802]<=16'd57308;
ROM1[2803]<=16'd4799; ROM2[2803]<=16'd0; ROM3[2803]<=16'd23824; ROM4[2803]<=16'd57318;
ROM1[2804]<=16'd4794; ROM2[2804]<=16'd0; ROM3[2804]<=16'd23841; ROM4[2804]<=16'd57327;
ROM1[2805]<=16'd4777; ROM2[2805]<=16'd0; ROM3[2805]<=16'd23832; ROM4[2805]<=16'd57315;
ROM1[2806]<=16'd4781; ROM2[2806]<=16'd0; ROM3[2806]<=16'd23820; ROM4[2806]<=16'd57307;
ROM1[2807]<=16'd4806; ROM2[2807]<=16'd0; ROM3[2807]<=16'd23796; ROM4[2807]<=16'd57299;
ROM1[2808]<=16'd4820; ROM2[2808]<=16'd0; ROM3[2808]<=16'd23783; ROM4[2808]<=16'd57294;
ROM1[2809]<=16'd4823; ROM2[2809]<=16'd0; ROM3[2809]<=16'd23795; ROM4[2809]<=16'd57304;
ROM1[2810]<=16'd4799; ROM2[2810]<=16'd0; ROM3[2810]<=16'd23800; ROM4[2810]<=16'd57306;
ROM1[2811]<=16'd4776; ROM2[2811]<=16'd0; ROM3[2811]<=16'd23805; ROM4[2811]<=16'd57303;
ROM1[2812]<=16'd4767; ROM2[2812]<=16'd0; ROM3[2812]<=16'd23814; ROM4[2812]<=16'd57309;
ROM1[2813]<=16'd4760; ROM2[2813]<=16'd0; ROM3[2813]<=16'd23819; ROM4[2813]<=16'd57310;
ROM1[2814]<=16'd4774; ROM2[2814]<=16'd0; ROM3[2814]<=16'd23824; ROM4[2814]<=16'd57314;
ROM1[2815]<=16'd4799; ROM2[2815]<=16'd0; ROM3[2815]<=16'd23812; ROM4[2815]<=16'd57314;
ROM1[2816]<=16'd4822; ROM2[2816]<=16'd0; ROM3[2816]<=16'd23793; ROM4[2816]<=16'd57308;
ROM1[2817]<=16'd4820; ROM2[2817]<=16'd0; ROM3[2817]<=16'd23790; ROM4[2817]<=16'd57308;
ROM1[2818]<=16'd4804; ROM2[2818]<=16'd0; ROM3[2818]<=16'd23800; ROM4[2818]<=16'd57307;
ROM1[2819]<=16'd4792; ROM2[2819]<=16'd0; ROM3[2819]<=16'd23814; ROM4[2819]<=16'd57316;
ROM1[2820]<=16'd4789; ROM2[2820]<=16'd0; ROM3[2820]<=16'd23827; ROM4[2820]<=16'd57326;
ROM1[2821]<=16'd4767; ROM2[2821]<=16'd0; ROM3[2821]<=16'd23819; ROM4[2821]<=16'd57314;
ROM1[2822]<=16'd4766; ROM2[2822]<=16'd0; ROM3[2822]<=16'd23810; ROM4[2822]<=16'd57307;
ROM1[2823]<=16'd4791; ROM2[2823]<=16'd0; ROM3[2823]<=16'd23806; ROM4[2823]<=16'd57307;
ROM1[2824]<=16'd4814; ROM2[2824]<=16'd0; ROM3[2824]<=16'd23792; ROM4[2824]<=16'd57303;
ROM1[2825]<=16'd4824; ROM2[2825]<=16'd0; ROM3[2825]<=16'd23792; ROM4[2825]<=16'd57307;
ROM1[2826]<=16'd4815; ROM2[2826]<=16'd0; ROM3[2826]<=16'd23799; ROM4[2826]<=16'd57312;
ROM1[2827]<=16'd4802; ROM2[2827]<=16'd0; ROM3[2827]<=16'd23807; ROM4[2827]<=16'd57310;
ROM1[2828]<=16'd4795; ROM2[2828]<=16'd0; ROM3[2828]<=16'd23816; ROM4[2828]<=16'd57308;
ROM1[2829]<=16'd4781; ROM2[2829]<=16'd0; ROM3[2829]<=16'd23823; ROM4[2829]<=16'd57310;
ROM1[2830]<=16'd4771; ROM2[2830]<=16'd0; ROM3[2830]<=16'd23816; ROM4[2830]<=16'd57309;
ROM1[2831]<=16'd4779; ROM2[2831]<=16'd0; ROM3[2831]<=16'd23801; ROM4[2831]<=16'd57298;
ROM1[2832]<=16'd4805; ROM2[2832]<=16'd0; ROM3[2832]<=16'd23779; ROM4[2832]<=16'd57288;
ROM1[2833]<=16'd4824; ROM2[2833]<=16'd0; ROM3[2833]<=16'd23771; ROM4[2833]<=16'd57292;
ROM1[2834]<=16'd4817; ROM2[2834]<=16'd0; ROM3[2834]<=16'd23783; ROM4[2834]<=16'd57295;
ROM1[2835]<=16'd4794; ROM2[2835]<=16'd0; ROM3[2835]<=16'd23787; ROM4[2835]<=16'd57294;
ROM1[2836]<=16'd4775; ROM2[2836]<=16'd0; ROM3[2836]<=16'd23792; ROM4[2836]<=16'd57292;
ROM1[2837]<=16'd4749; ROM2[2837]<=16'd0; ROM3[2837]<=16'd23787; ROM4[2837]<=16'd57274;
ROM1[2838]<=16'd4730; ROM2[2838]<=16'd0; ROM3[2838]<=16'd23778; ROM4[2838]<=16'd57263;
ROM1[2839]<=16'd4730; ROM2[2839]<=16'd0; ROM3[2839]<=16'd23770; ROM4[2839]<=16'd57255;
ROM1[2840]<=16'd4756; ROM2[2840]<=16'd0; ROM3[2840]<=16'd23757; ROM4[2840]<=16'd57249;
ROM1[2841]<=16'd4795; ROM2[2841]<=16'd0; ROM3[2841]<=16'd23757; ROM4[2841]<=16'd57261;
ROM1[2842]<=16'd4814; ROM2[2842]<=16'd0; ROM3[2842]<=16'd23771; ROM4[2842]<=16'd57274;
ROM1[2843]<=16'd4800; ROM2[2843]<=16'd0; ROM3[2843]<=16'd23781; ROM4[2843]<=16'd57278;
ROM1[2844]<=16'd4756; ROM2[2844]<=16'd0; ROM3[2844]<=16'd23772; ROM4[2844]<=16'd57261;
ROM1[2845]<=16'd4731; ROM2[2845]<=16'd0; ROM3[2845]<=16'd23770; ROM4[2845]<=16'd57251;
ROM1[2846]<=16'd4711; ROM2[2846]<=16'd0; ROM3[2846]<=16'd23769; ROM4[2846]<=16'd57245;
ROM1[2847]<=16'd4715; ROM2[2847]<=16'd0; ROM3[2847]<=16'd23765; ROM4[2847]<=16'd57241;
ROM1[2848]<=16'd4757; ROM2[2848]<=16'd0; ROM3[2848]<=16'd23775; ROM4[2848]<=16'd57256;
ROM1[2849]<=16'd4795; ROM2[2849]<=16'd0; ROM3[2849]<=16'd23772; ROM4[2849]<=16'd57264;
ROM1[2850]<=16'd4790; ROM2[2850]<=16'd0; ROM3[2850]<=16'd23750; ROM4[2850]<=16'd57253;
ROM1[2851]<=16'd4769; ROM2[2851]<=16'd0; ROM3[2851]<=16'd23747; ROM4[2851]<=16'd57249;
ROM1[2852]<=16'd4752; ROM2[2852]<=16'd0; ROM3[2852]<=16'd23756; ROM4[2852]<=16'd57252;
ROM1[2853]<=16'd4739; ROM2[2853]<=16'd0; ROM3[2853]<=16'd23760; ROM4[2853]<=16'd57248;
ROM1[2854]<=16'd4730; ROM2[2854]<=16'd0; ROM3[2854]<=16'd23776; ROM4[2854]<=16'd57259;
ROM1[2855]<=16'd4725; ROM2[2855]<=16'd0; ROM3[2855]<=16'd23786; ROM4[2855]<=16'd57266;
ROM1[2856]<=16'd4754; ROM2[2856]<=16'd0; ROM3[2856]<=16'd23793; ROM4[2856]<=16'd57277;
ROM1[2857]<=16'd4808; ROM2[2857]<=16'd0; ROM3[2857]<=16'd23800; ROM4[2857]<=16'd57301;
ROM1[2858]<=16'd4826; ROM2[2858]<=16'd0; ROM3[2858]<=16'd23790; ROM4[2858]<=16'd57297;
ROM1[2859]<=16'd4807; ROM2[2859]<=16'd0; ROM3[2859]<=16'd23784; ROM4[2859]<=16'd57289;
ROM1[2860]<=16'd4787; ROM2[2860]<=16'd0; ROM3[2860]<=16'd23787; ROM4[2860]<=16'd57285;
ROM1[2861]<=16'd4770; ROM2[2861]<=16'd0; ROM3[2861]<=16'd23791; ROM4[2861]<=16'd57282;
ROM1[2862]<=16'd4761; ROM2[2862]<=16'd0; ROM3[2862]<=16'd23803; ROM4[2862]<=16'd57287;
ROM1[2863]<=16'd4760; ROM2[2863]<=16'd0; ROM3[2863]<=16'd23812; ROM4[2863]<=16'd57290;
ROM1[2864]<=16'd4769; ROM2[2864]<=16'd0; ROM3[2864]<=16'd23810; ROM4[2864]<=16'd57291;
ROM1[2865]<=16'd4787; ROM2[2865]<=16'd0; ROM3[2865]<=16'd23792; ROM4[2865]<=16'd57283;
ROM1[2866]<=16'd4815; ROM2[2866]<=16'd0; ROM3[2866]<=16'd23787; ROM4[2866]<=16'd57287;
ROM1[2867]<=16'd4836; ROM2[2867]<=16'd0; ROM3[2867]<=16'd23809; ROM4[2867]<=16'd57309;
ROM1[2868]<=16'd4811; ROM2[2868]<=16'd0; ROM3[2868]<=16'd23811; ROM4[2868]<=16'd57303;
ROM1[2869]<=16'd4781; ROM2[2869]<=16'd0; ROM3[2869]<=16'd23804; ROM4[2869]<=16'd57291;
ROM1[2870]<=16'd4778; ROM2[2870]<=16'd0; ROM3[2870]<=16'd23817; ROM4[2870]<=16'd57297;
ROM1[2871]<=16'd4791; ROM2[2871]<=16'd0; ROM3[2871]<=16'd23848; ROM4[2871]<=16'd57320;
ROM1[2872]<=16'd4802; ROM2[2872]<=16'd0; ROM3[2872]<=16'd23854; ROM4[2872]<=16'd57330;
ROM1[2873]<=16'd4816; ROM2[2873]<=16'd0; ROM3[2873]<=16'd23839; ROM4[2873]<=16'd57323;
ROM1[2874]<=16'd4848; ROM2[2874]<=16'd0; ROM3[2874]<=16'd23826; ROM4[2874]<=16'd57324;
ROM1[2875]<=16'd4844; ROM2[2875]<=16'd0; ROM3[2875]<=16'd23810; ROM4[2875]<=16'd57315;
ROM1[2876]<=16'd4817; ROM2[2876]<=16'd0; ROM3[2876]<=16'd23801; ROM4[2876]<=16'd57301;
ROM1[2877]<=16'd4804; ROM2[2877]<=16'd0; ROM3[2877]<=16'd23808; ROM4[2877]<=16'd57299;
ROM1[2878]<=16'd4790; ROM2[2878]<=16'd0; ROM3[2878]<=16'd23816; ROM4[2878]<=16'd57303;
ROM1[2879]<=16'd4762; ROM2[2879]<=16'd0; ROM3[2879]<=16'd23811; ROM4[2879]<=16'd57292;
ROM1[2880]<=16'd4760; ROM2[2880]<=16'd0; ROM3[2880]<=16'd23812; ROM4[2880]<=16'd57292;
ROM1[2881]<=16'd4791; ROM2[2881]<=16'd0; ROM3[2881]<=16'd23818; ROM4[2881]<=16'd57308;
ROM1[2882]<=16'd4836; ROM2[2882]<=16'd0; ROM3[2882]<=16'd23810; ROM4[2882]<=16'd57312;
ROM1[2883]<=16'd4845; ROM2[2883]<=16'd0; ROM3[2883]<=16'd23785; ROM4[2883]<=16'd57297;
ROM1[2884]<=16'd4833; ROM2[2884]<=16'd0; ROM3[2884]<=16'd23787; ROM4[2884]<=16'd57301;
ROM1[2885]<=16'd4824; ROM2[2885]<=16'd0; ROM3[2885]<=16'd23803; ROM4[2885]<=16'd57310;
ROM1[2886]<=16'd4817; ROM2[2886]<=16'd0; ROM3[2886]<=16'd23813; ROM4[2886]<=16'd57314;
ROM1[2887]<=16'd4826; ROM2[2887]<=16'd0; ROM3[2887]<=16'd23839; ROM4[2887]<=16'd57330;
ROM1[2888]<=16'd4829; ROM2[2888]<=16'd0; ROM3[2888]<=16'd23857; ROM4[2888]<=16'd57341;
ROM1[2889]<=16'd4827; ROM2[2889]<=16'd0; ROM3[2889]<=16'd23847; ROM4[2889]<=16'd57332;
ROM1[2890]<=16'd4866; ROM2[2890]<=16'd0; ROM3[2890]<=16'd23826; ROM4[2890]<=16'd57323;
ROM1[2891]<=16'd4906; ROM2[2891]<=16'd0; ROM3[2891]<=16'd23807; ROM4[2891]<=16'd57322;
ROM1[2892]<=16'd4911; ROM2[2892]<=16'd0; ROM3[2892]<=16'd23802; ROM4[2892]<=16'd57318;
ROM1[2893]<=16'd4911; ROM2[2893]<=16'd0; ROM3[2893]<=16'd23819; ROM4[2893]<=16'd57326;
ROM1[2894]<=16'd4904; ROM2[2894]<=16'd0; ROM3[2894]<=16'd23837; ROM4[2894]<=16'd57332;
ROM1[2895]<=16'd4901; ROM2[2895]<=16'd0; ROM3[2895]<=16'd23847; ROM4[2895]<=16'd57337;
ROM1[2896]<=16'd4912; ROM2[2896]<=16'd0; ROM3[2896]<=16'd23865; ROM4[2896]<=16'd57351;
ROM1[2897]<=16'd4940; ROM2[2897]<=16'd0; ROM3[2897]<=16'd23869; ROM4[2897]<=16'd57363;
ROM1[2898]<=16'd4976; ROM2[2898]<=16'd0; ROM3[2898]<=16'd23859; ROM4[2898]<=16'd57368;
ROM1[2899]<=16'd5026; ROM2[2899]<=16'd0; ROM3[2899]<=16'd23845; ROM4[2899]<=16'd57369;
ROM1[2900]<=16'd5064; ROM2[2900]<=16'd0; ROM3[2900]<=16'd23844; ROM4[2900]<=16'd57376;
ROM1[2901]<=16'd5091; ROM2[2901]<=16'd0; ROM3[2901]<=16'd23870; ROM4[2901]<=16'd57400;
ROM1[2902]<=16'd5094; ROM2[2902]<=16'd0; ROM3[2902]<=16'd23888; ROM4[2902]<=16'd57415;
ROM1[2903]<=16'd5092; ROM2[2903]<=16'd0; ROM3[2903]<=16'd23892; ROM4[2903]<=16'd57414;
ROM1[2904]<=16'd5081; ROM2[2904]<=16'd0; ROM3[2904]<=16'd23885; ROM4[2904]<=16'd57405;
ROM1[2905]<=16'd5072; ROM2[2905]<=16'd0; ROM3[2905]<=16'd23864; ROM4[2905]<=16'd57389;
ROM1[2906]<=16'd5085; ROM2[2906]<=16'd0; ROM3[2906]<=16'd23844; ROM4[2906]<=16'd57376;
ROM1[2907]<=16'd5126; ROM2[2907]<=16'd0; ROM3[2907]<=16'd23828; ROM4[2907]<=16'd57375;
ROM1[2908]<=16'd5157; ROM2[2908]<=16'd0; ROM3[2908]<=16'd23825; ROM4[2908]<=16'd57376;
ROM1[2909]<=16'd5151; ROM2[2909]<=16'd0; ROM3[2909]<=16'd23826; ROM4[2909]<=16'd57371;
ROM1[2910]<=16'd5137; ROM2[2910]<=16'd0; ROM3[2910]<=16'd23831; ROM4[2910]<=16'd57374;
ROM1[2911]<=16'd5132; ROM2[2911]<=16'd0; ROM3[2911]<=16'd23837; ROM4[2911]<=16'd57375;
ROM1[2912]<=16'd5133; ROM2[2912]<=16'd0; ROM3[2912]<=16'd23838; ROM4[2912]<=16'd57377;
ROM1[2913]<=16'd5145; ROM2[2913]<=16'd0; ROM3[2913]<=16'd23847; ROM4[2913]<=16'd57387;
ROM1[2914]<=16'd5176; ROM2[2914]<=16'd0; ROM3[2914]<=16'd23855; ROM4[2914]<=16'd57398;
ROM1[2915]<=16'd5223; ROM2[2915]<=16'd0; ROM3[2915]<=16'd23854; ROM4[2915]<=16'd57410;
ROM1[2916]<=16'd5262; ROM2[2916]<=16'd0; ROM3[2916]<=16'd23850; ROM4[2916]<=16'd57415;
ROM1[2917]<=16'd5258; ROM2[2917]<=16'd0; ROM3[2917]<=16'd23841; ROM4[2917]<=16'd57407;
ROM1[2918]<=16'd5244; ROM2[2918]<=16'd0; ROM3[2918]<=16'd23847; ROM4[2918]<=16'd57405;
ROM1[2919]<=16'd5245; ROM2[2919]<=16'd0; ROM3[2919]<=16'd23864; ROM4[2919]<=16'd57413;
ROM1[2920]<=16'd5240; ROM2[2920]<=16'd0; ROM3[2920]<=16'd23861; ROM4[2920]<=16'd57407;
ROM1[2921]<=16'd5225; ROM2[2921]<=16'd0; ROM3[2921]<=16'd23853; ROM4[2921]<=16'd57393;
ROM1[2922]<=16'd5246; ROM2[2922]<=16'd0; ROM3[2922]<=16'd23856; ROM4[2922]<=16'd57398;
ROM1[2923]<=16'd5277; ROM2[2923]<=16'd0; ROM3[2923]<=16'd23848; ROM4[2923]<=16'd57405;
ROM1[2924]<=16'd5314; ROM2[2924]<=16'd0; ROM3[2924]<=16'd23837; ROM4[2924]<=16'd57411;
ROM1[2925]<=16'd5329; ROM2[2925]<=16'd0; ROM3[2925]<=16'd23837; ROM4[2925]<=16'd57418;
ROM1[2926]<=16'd5326; ROM2[2926]<=16'd0; ROM3[2926]<=16'd23838; ROM4[2926]<=16'd57421;
ROM1[2927]<=16'd5318; ROM2[2927]<=16'd0; ROM3[2927]<=16'd23846; ROM4[2927]<=16'd57423;
ROM1[2928]<=16'd5315; ROM2[2928]<=16'd0; ROM3[2928]<=16'd23862; ROM4[2928]<=16'd57435;
ROM1[2929]<=16'd5330; ROM2[2929]<=16'd0; ROM3[2929]<=16'd23891; ROM4[2929]<=16'd57460;
ROM1[2930]<=16'd5348; ROM2[2930]<=16'd0; ROM3[2930]<=16'd23906; ROM4[2930]<=16'd57472;
ROM1[2931]<=16'd5343; ROM2[2931]<=16'd0; ROM3[2931]<=16'd23880; ROM4[2931]<=16'd57456;
ROM1[2932]<=16'd5364; ROM2[2932]<=16'd0; ROM3[2932]<=16'd23858; ROM4[2932]<=16'd57441;
ROM1[2933]<=16'd5395; ROM2[2933]<=16'd0; ROM3[2933]<=16'd23860; ROM4[2933]<=16'd57450;
ROM1[2934]<=16'd5382; ROM2[2934]<=16'd0; ROM3[2934]<=16'd23862; ROM4[2934]<=16'd57450;
ROM1[2935]<=16'd5367; ROM2[2935]<=16'd0; ROM3[2935]<=16'd23874; ROM4[2935]<=16'd57451;
ROM1[2936]<=16'd5373; ROM2[2936]<=16'd0; ROM3[2936]<=16'd23902; ROM4[2936]<=16'd57472;
ROM1[2937]<=16'd5355; ROM2[2937]<=16'd0; ROM3[2937]<=16'd23908; ROM4[2937]<=16'd57470;
ROM1[2938]<=16'd5335; ROM2[2938]<=16'd0; ROM3[2938]<=16'd23900; ROM4[2938]<=16'd57458;
ROM1[2939]<=16'd5347; ROM2[2939]<=16'd0; ROM3[2939]<=16'd23903; ROM4[2939]<=16'd57462;
ROM1[2940]<=16'd5378; ROM2[2940]<=16'd0; ROM3[2940]<=16'd23896; ROM4[2940]<=16'd57465;
ROM1[2941]<=16'd5410; ROM2[2941]<=16'd0; ROM3[2941]<=16'd23887; ROM4[2941]<=16'd57467;
ROM1[2942]<=16'd5412; ROM2[2942]<=16'd0; ROM3[2942]<=16'd23894; ROM4[2942]<=16'd57472;
ROM1[2943]<=16'd5403; ROM2[2943]<=16'd0; ROM3[2943]<=16'd23912; ROM4[2943]<=16'd57483;
ROM1[2944]<=16'd5384; ROM2[2944]<=16'd0; ROM3[2944]<=16'd23919; ROM4[2944]<=16'd57483;
ROM1[2945]<=16'd5350; ROM2[2945]<=16'd0; ROM3[2945]<=16'd23910; ROM4[2945]<=16'd57468;
ROM1[2946]<=16'd5324; ROM2[2946]<=16'd0; ROM3[2946]<=16'd23903; ROM4[2946]<=16'd57459;
ROM1[2947]<=16'd5317; ROM2[2947]<=16'd0; ROM3[2947]<=16'd23895; ROM4[2947]<=16'd57454;
ROM1[2948]<=16'd5329; ROM2[2948]<=16'd0; ROM3[2948]<=16'd23886; ROM4[2948]<=16'd57450;
ROM1[2949]<=16'd5361; ROM2[2949]<=16'd0; ROM3[2949]<=16'd23875; ROM4[2949]<=16'd57453;
ROM1[2950]<=16'd5366; ROM2[2950]<=16'd0; ROM3[2950]<=16'd23871; ROM4[2950]<=16'd57450;
ROM1[2951]<=16'd5343; ROM2[2951]<=16'd0; ROM3[2951]<=16'd23873; ROM4[2951]<=16'd57441;
ROM1[2952]<=16'd5328; ROM2[2952]<=16'd0; ROM3[2952]<=16'd23886; ROM4[2952]<=16'd57445;
ROM1[2953]<=16'd5321; ROM2[2953]<=16'd0; ROM3[2953]<=16'd23901; ROM4[2953]<=16'd57459;
ROM1[2954]<=16'd5298; ROM2[2954]<=16'd0; ROM3[2954]<=16'd23908; ROM4[2954]<=16'd57463;
ROM1[2955]<=16'd5277; ROM2[2955]<=16'd0; ROM3[2955]<=16'd23902; ROM4[2955]<=16'd57455;
ROM1[2956]<=16'd5285; ROM2[2956]<=16'd0; ROM3[2956]<=16'd23887; ROM4[2956]<=16'd57445;
ROM1[2957]<=16'd5291; ROM2[2957]<=16'd0; ROM3[2957]<=16'd23863; ROM4[2957]<=16'd57427;
ROM1[2958]<=16'd5289; ROM2[2958]<=16'd0; ROM3[2958]<=16'd23849; ROM4[2958]<=16'd57415;
ROM1[2959]<=16'd5265; ROM2[2959]<=16'd0; ROM3[2959]<=16'd23850; ROM4[2959]<=16'd57413;
ROM1[2960]<=16'd5238; ROM2[2960]<=16'd0; ROM3[2960]<=16'd23856; ROM4[2960]<=16'd57411;
ROM1[2961]<=16'd5225; ROM2[2961]<=16'd0; ROM3[2961]<=16'd23877; ROM4[2961]<=16'd57423;
ROM1[2962]<=16'd5193; ROM2[2962]<=16'd0; ROM3[2962]<=16'd23874; ROM4[2962]<=16'd57418;
ROM1[2963]<=16'd5175; ROM2[2963]<=16'd0; ROM3[2963]<=16'd23875; ROM4[2963]<=16'd57413;
ROM1[2964]<=16'd5176; ROM2[2964]<=16'd0; ROM3[2964]<=16'd23878; ROM4[2964]<=16'd57417;
ROM1[2965]<=16'd5169; ROM2[2965]<=16'd0; ROM3[2965]<=16'd23839; ROM4[2965]<=16'd57390;
ROM1[2966]<=16'd5181; ROM2[2966]<=16'd0; ROM3[2966]<=16'd23816; ROM4[2966]<=16'd57376;
ROM1[2967]<=16'd5184; ROM2[2967]<=16'd0; ROM3[2967]<=16'd23826; ROM4[2967]<=16'd57390;
ROM1[2968]<=16'd5158; ROM2[2968]<=16'd0; ROM3[2968]<=16'd23833; ROM4[2968]<=16'd57393;
ROM1[2969]<=16'd5133; ROM2[2969]<=16'd0; ROM3[2969]<=16'd23841; ROM4[2969]<=16'd57394;
ROM1[2970]<=16'd5121; ROM2[2970]<=16'd0; ROM3[2970]<=16'd23857; ROM4[2970]<=16'd57403;
ROM1[2971]<=16'd5095; ROM2[2971]<=16'd0; ROM3[2971]<=16'd23861; ROM4[2971]<=16'd57398;
ROM1[2972]<=16'd5085; ROM2[2972]<=16'd0; ROM3[2972]<=16'd23853; ROM4[2972]<=16'd57391;
ROM1[2973]<=16'd5102; ROM2[2973]<=16'd0; ROM3[2973]<=16'd23844; ROM4[2973]<=16'd57388;
ROM1[2974]<=16'd5120; ROM2[2974]<=16'd0; ROM3[2974]<=16'd23828; ROM4[2974]<=16'd57378;
ROM1[2975]<=16'd5110; ROM2[2975]<=16'd0; ROM3[2975]<=16'd23814; ROM4[2975]<=16'd57368;
ROM1[2976]<=16'd5081; ROM2[2976]<=16'd0; ROM3[2976]<=16'd23815; ROM4[2976]<=16'd57362;
ROM1[2977]<=16'd5060; ROM2[2977]<=16'd0; ROM3[2977]<=16'd23830; ROM4[2977]<=16'd57366;
ROM1[2978]<=16'd5056; ROM2[2978]<=16'd0; ROM3[2978]<=16'd23853; ROM4[2978]<=16'd57385;
ROM1[2979]<=16'd5048; ROM2[2979]<=16'd0; ROM3[2979]<=16'd23872; ROM4[2979]<=16'd57394;
ROM1[2980]<=16'd5020; ROM2[2980]<=16'd0; ROM3[2980]<=16'd23851; ROM4[2980]<=16'd57371;
ROM1[2981]<=16'd5022; ROM2[2981]<=16'd0; ROM3[2981]<=16'd23831; ROM4[2981]<=16'd57359;
ROM1[2982]<=16'd5048; ROM2[2982]<=16'd0; ROM3[2982]<=16'd23817; ROM4[2982]<=16'd57354;
ROM1[2983]<=16'd5048; ROM2[2983]<=16'd0; ROM3[2983]<=16'd23794; ROM4[2983]<=16'd57340;
ROM1[2984]<=16'd5035; ROM2[2984]<=16'd0; ROM3[2984]<=16'd23800; ROM4[2984]<=16'd57346;
ROM1[2985]<=16'd5015; ROM2[2985]<=16'd0; ROM3[2985]<=16'd23814; ROM4[2985]<=16'd57350;
ROM1[2986]<=16'd4993; ROM2[2986]<=16'd0; ROM3[2986]<=16'd23817; ROM4[2986]<=16'd57346;
ROM1[2987]<=16'd4975; ROM2[2987]<=16'd0; ROM3[2987]<=16'd23827; ROM4[2987]<=16'd57351;
ROM1[2988]<=16'd4968; ROM2[2988]<=16'd0; ROM3[2988]<=16'd23837; ROM4[2988]<=16'd57356;
ROM1[2989]<=16'd4986; ROM2[2989]<=16'd0; ROM3[2989]<=16'd23845; ROM4[2989]<=16'd57365;
ROM1[2990]<=16'd5014; ROM2[2990]<=16'd0; ROM3[2990]<=16'd23841; ROM4[2990]<=16'd57369;
ROM1[2991]<=16'd5040; ROM2[2991]<=16'd0; ROM3[2991]<=16'd23830; ROM4[2991]<=16'd57367;
ROM1[2992]<=16'd5049; ROM2[2992]<=16'd0; ROM3[2992]<=16'd23847; ROM4[2992]<=16'd57380;
ROM1[2993]<=16'd5012; ROM2[2993]<=16'd0; ROM3[2993]<=16'd23845; ROM4[2993]<=16'd57371;
ROM1[2994]<=16'd4980; ROM2[2994]<=16'd0; ROM3[2994]<=16'd23842; ROM4[2994]<=16'd57364;
ROM1[2995]<=16'd4969; ROM2[2995]<=16'd0; ROM3[2995]<=16'd23849; ROM4[2995]<=16'd57366;
ROM1[2996]<=16'd4941; ROM2[2996]<=16'd0; ROM3[2996]<=16'd23839; ROM4[2996]<=16'd57347;
ROM1[2997]<=16'd4941; ROM2[2997]<=16'd0; ROM3[2997]<=16'd23835; ROM4[2997]<=16'd57345;
ROM1[2998]<=16'd4974; ROM2[2998]<=16'd0; ROM3[2998]<=16'd23836; ROM4[2998]<=16'd57347;
ROM1[2999]<=16'd5011; ROM2[2999]<=16'd0; ROM3[2999]<=16'd23832; ROM4[2999]<=16'd57353;
ROM1[3000]<=16'd5012; ROM2[3000]<=16'd0; ROM3[3000]<=16'd23826; ROM4[3000]<=16'd57350;
ROM1[3001]<=16'd4986; ROM2[3001]<=16'd0; ROM3[3001]<=16'd23817; ROM4[3001]<=16'd57337;
ROM1[3002]<=16'd4962; ROM2[3002]<=16'd0; ROM3[3002]<=16'd23817; ROM4[3002]<=16'd57334;
ROM1[3003]<=16'd4949; ROM2[3003]<=16'd0; ROM3[3003]<=16'd23826; ROM4[3003]<=16'd57336;
ROM1[3004]<=16'd4945; ROM2[3004]<=16'd0; ROM3[3004]<=16'd23840; ROM4[3004]<=16'd57349;
ROM1[3005]<=16'd4950; ROM2[3005]<=16'd0; ROM3[3005]<=16'd23857; ROM4[3005]<=16'd57357;
ROM1[3006]<=16'd4950; ROM2[3006]<=16'd0; ROM3[3006]<=16'd23840; ROM4[3006]<=16'd57343;
ROM1[3007]<=16'd4959; ROM2[3007]<=16'd0; ROM3[3007]<=16'd23807; ROM4[3007]<=16'd57323;
ROM1[3008]<=16'd4955; ROM2[3008]<=16'd0; ROM3[3008]<=16'd23780; ROM4[3008]<=16'd57299;
ROM1[3009]<=16'd4925; ROM2[3009]<=16'd0; ROM3[3009]<=16'd23768; ROM4[3009]<=16'd57284;
ROM1[3010]<=16'd4904; ROM2[3010]<=16'd0; ROM3[3010]<=16'd23768; ROM4[3010]<=16'd57278;
ROM1[3011]<=16'd4886; ROM2[3011]<=16'd0; ROM3[3011]<=16'd23767; ROM4[3011]<=16'd57270;
ROM1[3012]<=16'd4863; ROM2[3012]<=16'd0; ROM3[3012]<=16'd23769; ROM4[3012]<=16'd57267;
ROM1[3013]<=16'd4859; ROM2[3013]<=16'd0; ROM3[3013]<=16'd23776; ROM4[3013]<=16'd57273;
ROM1[3014]<=16'd4880; ROM2[3014]<=16'd0; ROM3[3014]<=16'd23784; ROM4[3014]<=16'd57284;
ROM1[3015]<=16'd4896; ROM2[3015]<=16'd0; ROM3[3015]<=16'd23767; ROM4[3015]<=16'd57274;
ROM1[3016]<=16'd4906; ROM2[3016]<=16'd0; ROM3[3016]<=16'd23748; ROM4[3016]<=16'd57262;
ROM1[3017]<=16'd4906; ROM2[3017]<=16'd0; ROM3[3017]<=16'd23757; ROM4[3017]<=16'd57271;
ROM1[3018]<=16'd4891; ROM2[3018]<=16'd0; ROM3[3018]<=16'd23772; ROM4[3018]<=16'd57284;
ROM1[3019]<=16'd4883; ROM2[3019]<=16'd0; ROM3[3019]<=16'd23791; ROM4[3019]<=16'd57296;
ROM1[3020]<=16'd4874; ROM2[3020]<=16'd0; ROM3[3020]<=16'd23797; ROM4[3020]<=16'd57298;
ROM1[3021]<=16'd4862; ROM2[3021]<=16'd0; ROM3[3021]<=16'd23804; ROM4[3021]<=16'd57298;
ROM1[3022]<=16'd4877; ROM2[3022]<=16'd0; ROM3[3022]<=16'd23820; ROM4[3022]<=16'd57311;
ROM1[3023]<=16'd4895; ROM2[3023]<=16'd0; ROM3[3023]<=16'd23813; ROM4[3023]<=16'd57312;
ROM1[3024]<=16'd4927; ROM2[3024]<=16'd0; ROM3[3024]<=16'd23806; ROM4[3024]<=16'd57316;
ROM1[3025]<=16'd4932; ROM2[3025]<=16'd0; ROM3[3025]<=16'd23799; ROM4[3025]<=16'd57316;
ROM1[3026]<=16'd4902; ROM2[3026]<=16'd0; ROM3[3026]<=16'd23789; ROM4[3026]<=16'd57301;
ROM1[3027]<=16'd4878; ROM2[3027]<=16'd0; ROM3[3027]<=16'd23794; ROM4[3027]<=16'd57296;
ROM1[3028]<=16'd4868; ROM2[3028]<=16'd0; ROM3[3028]<=16'd23801; ROM4[3028]<=16'd57299;
ROM1[3029]<=16'd4852; ROM2[3029]<=16'd0; ROM3[3029]<=16'd23804; ROM4[3029]<=16'd57293;
ROM1[3030]<=16'd4838; ROM2[3030]<=16'd0; ROM3[3030]<=16'd23794; ROM4[3030]<=16'd57284;
ROM1[3031]<=16'd4856; ROM2[3031]<=16'd0; ROM3[3031]<=16'd23789; ROM4[3031]<=16'd57283;
ROM1[3032]<=16'd4891; ROM2[3032]<=16'd0; ROM3[3032]<=16'd23786; ROM4[3032]<=16'd57288;
ROM1[3033]<=16'd4905; ROM2[3033]<=16'd0; ROM3[3033]<=16'd23777; ROM4[3033]<=16'd57290;
ROM1[3034]<=16'd4900; ROM2[3034]<=16'd0; ROM3[3034]<=16'd23787; ROM4[3034]<=16'd57293;
ROM1[3035]<=16'd4890; ROM2[3035]<=16'd0; ROM3[3035]<=16'd23809; ROM4[3035]<=16'd57304;
ROM1[3036]<=16'd4886; ROM2[3036]<=16'd0; ROM3[3036]<=16'd23826; ROM4[3036]<=16'd57313;
ROM1[3037]<=16'd4875; ROM2[3037]<=16'd0; ROM3[3037]<=16'd23837; ROM4[3037]<=16'd57313;
ROM1[3038]<=16'd4871; ROM2[3038]<=16'd0; ROM3[3038]<=16'd23844; ROM4[3038]<=16'd57320;
ROM1[3039]<=16'd4888; ROM2[3039]<=16'd0; ROM3[3039]<=16'd23847; ROM4[3039]<=16'd57330;
ROM1[3040]<=16'd4918; ROM2[3040]<=16'd0; ROM3[3040]<=16'd23840; ROM4[3040]<=16'd57331;
ROM1[3041]<=16'd4935; ROM2[3041]<=16'd0; ROM3[3041]<=16'd23820; ROM4[3041]<=16'd57320;
ROM1[3042]<=16'd4919; ROM2[3042]<=16'd0; ROM3[3042]<=16'd23810; ROM4[3042]<=16'd57307;
ROM1[3043]<=16'd4893; ROM2[3043]<=16'd0; ROM3[3043]<=16'd23809; ROM4[3043]<=16'd57301;
ROM1[3044]<=16'd4885; ROM2[3044]<=16'd0; ROM3[3044]<=16'd23821; ROM4[3044]<=16'd57307;
ROM1[3045]<=16'd4900; ROM2[3045]<=16'd0; ROM3[3045]<=16'd23853; ROM4[3045]<=16'd57339;
ROM1[3046]<=16'd4909; ROM2[3046]<=16'd0; ROM3[3046]<=16'd23879; ROM4[3046]<=16'd57359;
ROM1[3047]<=16'd4889; ROM2[3047]<=16'd0; ROM3[3047]<=16'd23856; ROM4[3047]<=16'd57336;
ROM1[3048]<=16'd4877; ROM2[3048]<=16'd0; ROM3[3048]<=16'd23818; ROM4[3048]<=16'd57305;
ROM1[3049]<=16'd4904; ROM2[3049]<=16'd0; ROM3[3049]<=16'd23808; ROM4[3049]<=16'd57305;
ROM1[3050]<=16'd4900; ROM2[3050]<=16'd0; ROM3[3050]<=16'd23806; ROM4[3050]<=16'd57305;
ROM1[3051]<=16'd4886; ROM2[3051]<=16'd0; ROM3[3051]<=16'd23813; ROM4[3051]<=16'd57313;
ROM1[3052]<=16'd4879; ROM2[3052]<=16'd0; ROM3[3052]<=16'd23828; ROM4[3052]<=16'd57324;
ROM1[3053]<=16'd4848; ROM2[3053]<=16'd0; ROM3[3053]<=16'd23820; ROM4[3053]<=16'd57316;
ROM1[3054]<=16'd4819; ROM2[3054]<=16'd0; ROM3[3054]<=16'd23814; ROM4[3054]<=16'd57310;
ROM1[3055]<=16'd4827; ROM2[3055]<=16'd0; ROM3[3055]<=16'd23830; ROM4[3055]<=16'd57321;
ROM1[3056]<=16'd4853; ROM2[3056]<=16'd0; ROM3[3056]<=16'd23839; ROM4[3056]<=16'd57335;
ROM1[3057]<=16'd4852; ROM2[3057]<=16'd0; ROM3[3057]<=16'd23794; ROM4[3057]<=16'd57304;
ROM1[3058]<=16'd4847; ROM2[3058]<=16'd0; ROM3[3058]<=16'd23759; ROM4[3058]<=16'd57278;
ROM1[3059]<=16'd4839; ROM2[3059]<=16'd0; ROM3[3059]<=16'd23757; ROM4[3059]<=16'd57274;
ROM1[3060]<=16'd4815; ROM2[3060]<=16'd0; ROM3[3060]<=16'd23758; ROM4[3060]<=16'd57270;
ROM1[3061]<=16'd4808; ROM2[3061]<=16'd0; ROM3[3061]<=16'd23775; ROM4[3061]<=16'd57277;
ROM1[3062]<=16'd4816; ROM2[3062]<=16'd0; ROM3[3062]<=16'd23796; ROM4[3062]<=16'd57291;
ROM1[3063]<=16'd4815; ROM2[3063]<=16'd0; ROM3[3063]<=16'd23809; ROM4[3063]<=16'd57298;
ROM1[3064]<=16'd4811; ROM2[3064]<=16'd0; ROM3[3064]<=16'd23793; ROM4[3064]<=16'd57282;
ROM1[3065]<=16'd4844; ROM2[3065]<=16'd0; ROM3[3065]<=16'd23781; ROM4[3065]<=16'd57279;
ROM1[3066]<=16'd4881; ROM2[3066]<=16'd0; ROM3[3066]<=16'd23780; ROM4[3066]<=16'd57286;
ROM1[3067]<=16'd4866; ROM2[3067]<=16'd0; ROM3[3067]<=16'd23767; ROM4[3067]<=16'd57269;
ROM1[3068]<=16'd4848; ROM2[3068]<=16'd0; ROM3[3068]<=16'd23773; ROM4[3068]<=16'd57267;
ROM1[3069]<=16'd4841; ROM2[3069]<=16'd0; ROM3[3069]<=16'd23791; ROM4[3069]<=16'd57275;
ROM1[3070]<=16'd4821; ROM2[3070]<=16'd0; ROM3[3070]<=16'd23792; ROM4[3070]<=16'd57267;
ROM1[3071]<=16'd4813; ROM2[3071]<=16'd0; ROM3[3071]<=16'd23800; ROM4[3071]<=16'd57271;
ROM1[3072]<=16'd4824; ROM2[3072]<=16'd0; ROM3[3072]<=16'd23805; ROM4[3072]<=16'd57277;
ROM1[3073]<=16'd4850; ROM2[3073]<=16'd0; ROM3[3073]<=16'd23805; ROM4[3073]<=16'd57282;
ROM1[3074]<=16'd4875; ROM2[3074]<=16'd0; ROM3[3074]<=16'd23798; ROM4[3074]<=16'd57282;
ROM1[3075]<=16'd4862; ROM2[3075]<=16'd0; ROM3[3075]<=16'd23784; ROM4[3075]<=16'd57265;
ROM1[3076]<=16'd4849; ROM2[3076]<=16'd0; ROM3[3076]<=16'd23796; ROM4[3076]<=16'd57268;
ROM1[3077]<=16'd4834; ROM2[3077]<=16'd0; ROM3[3077]<=16'd23809; ROM4[3077]<=16'd57270;
ROM1[3078]<=16'd4812; ROM2[3078]<=16'd0; ROM3[3078]<=16'd23810; ROM4[3078]<=16'd57260;
ROM1[3079]<=16'd4788; ROM2[3079]<=16'd0; ROM3[3079]<=16'd23808; ROM4[3079]<=16'd57250;
ROM1[3080]<=16'd4775; ROM2[3080]<=16'd0; ROM3[3080]<=16'd23800; ROM4[3080]<=16'd57240;
ROM1[3081]<=16'd4793; ROM2[3081]<=16'd0; ROM3[3081]<=16'd23795; ROM4[3081]<=16'd57240;
ROM1[3082]<=16'd4840; ROM2[3082]<=16'd0; ROM3[3082]<=16'd23792; ROM4[3082]<=16'd57253;
ROM1[3083]<=16'd4867; ROM2[3083]<=16'd0; ROM3[3083]<=16'd23792; ROM4[3083]<=16'd57265;
ROM1[3084]<=16'd4826; ROM2[3084]<=16'd0; ROM3[3084]<=16'd23769; ROM4[3084]<=16'd57242;
ROM1[3085]<=16'd4791; ROM2[3085]<=16'd0; ROM3[3085]<=16'd23760; ROM4[3085]<=16'd57227;
ROM1[3086]<=16'd4786; ROM2[3086]<=16'd0; ROM3[3086]<=16'd23776; ROM4[3086]<=16'd57236;
ROM1[3087]<=16'd4781; ROM2[3087]<=16'd0; ROM3[3087]<=16'd23796; ROM4[3087]<=16'd57254;
ROM1[3088]<=16'd4796; ROM2[3088]<=16'd0; ROM3[3088]<=16'd23822; ROM4[3088]<=16'd57282;
ROM1[3089]<=16'd4821; ROM2[3089]<=16'd0; ROM3[3089]<=16'd23835; ROM4[3089]<=16'd57298;
ROM1[3090]<=16'd4842; ROM2[3090]<=16'd0; ROM3[3090]<=16'd23824; ROM4[3090]<=16'd57299;
ROM1[3091]<=16'd4869; ROM2[3091]<=16'd0; ROM3[3091]<=16'd23819; ROM4[3091]<=16'd57308;
ROM1[3092]<=16'd4878; ROM2[3092]<=16'd0; ROM3[3092]<=16'd23830; ROM4[3092]<=16'd57323;
ROM1[3093]<=16'd4874; ROM2[3093]<=16'd0; ROM3[3093]<=16'd23848; ROM4[3093]<=16'd57340;
ROM1[3094]<=16'd4857; ROM2[3094]<=16'd0; ROM3[3094]<=16'd23855; ROM4[3094]<=16'd57340;
ROM1[3095]<=16'd4835; ROM2[3095]<=16'd0; ROM3[3095]<=16'd23851; ROM4[3095]<=16'd57331;
ROM1[3096]<=16'd4829; ROM2[3096]<=16'd0; ROM3[3096]<=16'd23859; ROM4[3096]<=16'd57336;
ROM1[3097]<=16'd4834; ROM2[3097]<=16'd0; ROM3[3097]<=16'd23859; ROM4[3097]<=16'd57338;
ROM1[3098]<=16'd4865; ROM2[3098]<=16'd0; ROM3[3098]<=16'd23850; ROM4[3098]<=16'd57344;
ROM1[3099]<=16'd4900; ROM2[3099]<=16'd0; ROM3[3099]<=16'd23836; ROM4[3099]<=16'd57342;
ROM1[3100]<=16'd4899; ROM2[3100]<=16'd0; ROM3[3100]<=16'd23826; ROM4[3100]<=16'd57333;
ROM1[3101]<=16'd4880; ROM2[3101]<=16'd0; ROM3[3101]<=16'd23827; ROM4[3101]<=16'd57331;
ROM1[3102]<=16'd4854; ROM2[3102]<=16'd0; ROM3[3102]<=16'd23828; ROM4[3102]<=16'd57323;
ROM1[3103]<=16'd4850; ROM2[3103]<=16'd0; ROM3[3103]<=16'd23838; ROM4[3103]<=16'd57329;
ROM1[3104]<=16'd4850; ROM2[3104]<=16'd0; ROM3[3104]<=16'd23848; ROM4[3104]<=16'd57339;
ROM1[3105]<=16'd4845; ROM2[3105]<=16'd0; ROM3[3105]<=16'd23847; ROM4[3105]<=16'd57332;
ROM1[3106]<=16'd4855; ROM2[3106]<=16'd0; ROM3[3106]<=16'd23833; ROM4[3106]<=16'd57326;
ROM1[3107]<=16'd4877; ROM2[3107]<=16'd0; ROM3[3107]<=16'd23806; ROM4[3107]<=16'd57315;
ROM1[3108]<=16'd4880; ROM2[3108]<=16'd0; ROM3[3108]<=16'd23786; ROM4[3108]<=16'd57297;
ROM1[3109]<=16'd4856; ROM2[3109]<=16'd0; ROM3[3109]<=16'd23778; ROM4[3109]<=16'd57288;
ROM1[3110]<=16'd4836; ROM2[3110]<=16'd0; ROM3[3110]<=16'd23784; ROM4[3110]<=16'd57285;
ROM1[3111]<=16'd4830; ROM2[3111]<=16'd0; ROM3[3111]<=16'd23802; ROM4[3111]<=16'd57291;
ROM1[3112]<=16'd4816; ROM2[3112]<=16'd0; ROM3[3112]<=16'd23810; ROM4[3112]<=16'd57293;
ROM1[3113]<=16'd4802; ROM2[3113]<=16'd0; ROM3[3113]<=16'd23806; ROM4[3113]<=16'd57286;
ROM1[3114]<=16'd4809; ROM2[3114]<=16'd0; ROM3[3114]<=16'd23800; ROM4[3114]<=16'd57278;
ROM1[3115]<=16'd4834; ROM2[3115]<=16'd0; ROM3[3115]<=16'd23787; ROM4[3115]<=16'd57272;
ROM1[3116]<=16'd4866; ROM2[3116]<=16'd0; ROM3[3116]<=16'd23782; ROM4[3116]<=16'd57276;
ROM1[3117]<=16'd4873; ROM2[3117]<=16'd0; ROM3[3117]<=16'd23790; ROM4[3117]<=16'd57282;
ROM1[3118]<=16'd4845; ROM2[3118]<=16'd0; ROM3[3118]<=16'd23785; ROM4[3118]<=16'd57274;
ROM1[3119]<=16'd4813; ROM2[3119]<=16'd0; ROM3[3119]<=16'd23778; ROM4[3119]<=16'd57263;
ROM1[3120]<=16'd4816; ROM2[3120]<=16'd0; ROM3[3120]<=16'd23799; ROM4[3120]<=16'd57277;
ROM1[3121]<=16'd4806; ROM2[3121]<=16'd0; ROM3[3121]<=16'd23803; ROM4[3121]<=16'd57279;
ROM1[3122]<=16'd4793; ROM2[3122]<=16'd0; ROM3[3122]<=16'd23791; ROM4[3122]<=16'd57266;
ROM1[3123]<=16'd4809; ROM2[3123]<=16'd0; ROM3[3123]<=16'd23778; ROM4[3123]<=16'd57260;
ROM1[3124]<=16'd4839; ROM2[3124]<=16'd0; ROM3[3124]<=16'd23766; ROM4[3124]<=16'd57262;
ROM1[3125]<=16'd4847; ROM2[3125]<=16'd0; ROM3[3125]<=16'd23764; ROM4[3125]<=16'd57263;
ROM1[3126]<=16'd4838; ROM2[3126]<=16'd0; ROM3[3126]<=16'd23775; ROM4[3126]<=16'd57267;
ROM1[3127]<=16'd4830; ROM2[3127]<=16'd0; ROM3[3127]<=16'd23793; ROM4[3127]<=16'd57278;
ROM1[3128]<=16'd4810; ROM2[3128]<=16'd0; ROM3[3128]<=16'd23792; ROM4[3128]<=16'd57274;
ROM1[3129]<=16'd4799; ROM2[3129]<=16'd0; ROM3[3129]<=16'd23798; ROM4[3129]<=16'd57275;
ROM1[3130]<=16'd4810; ROM2[3130]<=16'd0; ROM3[3130]<=16'd23810; ROM4[3130]<=16'd57292;
ROM1[3131]<=16'd4835; ROM2[3131]<=16'd0; ROM3[3131]<=16'd23812; ROM4[3131]<=16'd57301;
ROM1[3132]<=16'd4867; ROM2[3132]<=16'd0; ROM3[3132]<=16'd23801; ROM4[3132]<=16'd57301;
ROM1[3133]<=16'd4898; ROM2[3133]<=16'd0; ROM3[3133]<=16'd23814; ROM4[3133]<=16'd57320;
ROM1[3134]<=16'd4900; ROM2[3134]<=16'd0; ROM3[3134]<=16'd23833; ROM4[3134]<=16'd57337;
ROM1[3135]<=16'd4881; ROM2[3135]<=16'd0; ROM3[3135]<=16'd23840; ROM4[3135]<=16'd57342;
ROM1[3136]<=16'd4864; ROM2[3136]<=16'd0; ROM3[3136]<=16'd23841; ROM4[3136]<=16'd57337;
ROM1[3137]<=16'd4841; ROM2[3137]<=16'd0; ROM3[3137]<=16'd23839; ROM4[3137]<=16'd57331;
ROM1[3138]<=16'd4829; ROM2[3138]<=16'd0; ROM3[3138]<=16'd23842; ROM4[3138]<=16'd57332;
ROM1[3139]<=16'd4842; ROM2[3139]<=16'd0; ROM3[3139]<=16'd23843; ROM4[3139]<=16'd57337;
ROM1[3140]<=16'd4886; ROM2[3140]<=16'd0; ROM3[3140]<=16'd23851; ROM4[3140]<=16'd57354;
ROM1[3141]<=16'd4912; ROM2[3141]<=16'd0; ROM3[3141]<=16'd23833; ROM4[3141]<=16'd57352;
ROM1[3142]<=16'd4889; ROM2[3142]<=16'd0; ROM3[3142]<=16'd23809; ROM4[3142]<=16'd57330;
ROM1[3143]<=16'd4867; ROM2[3143]<=16'd0; ROM3[3143]<=16'd23814; ROM4[3143]<=16'd57325;
ROM1[3144]<=16'd4843; ROM2[3144]<=16'd0; ROM3[3144]<=16'd23816; ROM4[3144]<=16'd57320;
ROM1[3145]<=16'd4819; ROM2[3145]<=16'd0; ROM3[3145]<=16'd23815; ROM4[3145]<=16'd57312;
ROM1[3146]<=16'd4812; ROM2[3146]<=16'd0; ROM3[3146]<=16'd23825; ROM4[3146]<=16'd57313;
ROM1[3147]<=16'd4821; ROM2[3147]<=16'd0; ROM3[3147]<=16'd23830; ROM4[3147]<=16'd57314;
ROM1[3148]<=16'd4838; ROM2[3148]<=16'd0; ROM3[3148]<=16'd23819; ROM4[3148]<=16'd57306;
ROM1[3149]<=16'd4864; ROM2[3149]<=16'd0; ROM3[3149]<=16'd23805; ROM4[3149]<=16'd57302;
ROM1[3150]<=16'd4864; ROM2[3150]<=16'd0; ROM3[3150]<=16'd23796; ROM4[3150]<=16'd57297;
ROM1[3151]<=16'd4847; ROM2[3151]<=16'd0; ROM3[3151]<=16'd23797; ROM4[3151]<=16'd57293;
ROM1[3152]<=16'd4827; ROM2[3152]<=16'd0; ROM3[3152]<=16'd23805; ROM4[3152]<=16'd57288;
ROM1[3153]<=16'd4792; ROM2[3153]<=16'd0; ROM3[3153]<=16'd23788; ROM4[3153]<=16'd57261;
ROM1[3154]<=16'd4776; ROM2[3154]<=16'd0; ROM3[3154]<=16'd23785; ROM4[3154]<=16'd57257;
ROM1[3155]<=16'd4777; ROM2[3155]<=16'd0; ROM3[3155]<=16'd23786; ROM4[3155]<=16'd57259;
ROM1[3156]<=16'd4786; ROM2[3156]<=16'd0; ROM3[3156]<=16'd23767; ROM4[3156]<=16'd57250;
ROM1[3157]<=16'd4831; ROM2[3157]<=16'd0; ROM3[3157]<=16'd23762; ROM4[3157]<=16'd57261;
ROM1[3158]<=16'd4868; ROM2[3158]<=16'd0; ROM3[3158]<=16'd23772; ROM4[3158]<=16'd57279;
ROM1[3159]<=16'd4858; ROM2[3159]<=16'd0; ROM3[3159]<=16'd23780; ROM4[3159]<=16'd57284;
ROM1[3160]<=16'd4819; ROM2[3160]<=16'd0; ROM3[3160]<=16'd23771; ROM4[3160]<=16'd57267;
ROM1[3161]<=16'd4804; ROM2[3161]<=16'd0; ROM3[3161]<=16'd23779; ROM4[3161]<=16'd57268;
ROM1[3162]<=16'd4791; ROM2[3162]<=16'd0; ROM3[3162]<=16'd23789; ROM4[3162]<=16'd57273;
ROM1[3163]<=16'd4788; ROM2[3163]<=16'd0; ROM3[3163]<=16'd23792; ROM4[3163]<=16'd57274;
ROM1[3164]<=16'd4816; ROM2[3164]<=16'd0; ROM3[3164]<=16'd23797; ROM4[3164]<=16'd57284;
ROM1[3165]<=16'd4854; ROM2[3165]<=16'd0; ROM3[3165]<=16'd23794; ROM4[3165]<=16'd57290;
ROM1[3166]<=16'd4884; ROM2[3166]<=16'd0; ROM3[3166]<=16'd23788; ROM4[3166]<=16'd57295;
ROM1[3167]<=16'd4882; ROM2[3167]<=16'd0; ROM3[3167]<=16'd23789; ROM4[3167]<=16'd57298;
ROM1[3168]<=16'd4867; ROM2[3168]<=16'd0; ROM3[3168]<=16'd23797; ROM4[3168]<=16'd57297;
ROM1[3169]<=16'd4846; ROM2[3169]<=16'd0; ROM3[3169]<=16'd23801; ROM4[3169]<=16'd57289;
ROM1[3170]<=16'd4829; ROM2[3170]<=16'd0; ROM3[3170]<=16'd23801; ROM4[3170]<=16'd57284;
ROM1[3171]<=16'd4816; ROM2[3171]<=16'd0; ROM3[3171]<=16'd23805; ROM4[3171]<=16'd57279;
ROM1[3172]<=16'd4824; ROM2[3172]<=16'd0; ROM3[3172]<=16'd23806; ROM4[3172]<=16'd57285;
ROM1[3173]<=16'd4864; ROM2[3173]<=16'd0; ROM3[3173]<=16'd23813; ROM4[3173]<=16'd57306;
ROM1[3174]<=16'd4895; ROM2[3174]<=16'd0; ROM3[3174]<=16'd23801; ROM4[3174]<=16'd57306;
ROM1[3175]<=16'd4881; ROM2[3175]<=16'd0; ROM3[3175]<=16'd23781; ROM4[3175]<=16'd57291;
ROM1[3176]<=16'd4868; ROM2[3176]<=16'd0; ROM3[3176]<=16'd23791; ROM4[3176]<=16'd57293;
ROM1[3177]<=16'd4856; ROM2[3177]<=16'd0; ROM3[3177]<=16'd23804; ROM4[3177]<=16'd57297;
ROM1[3178]<=16'd4836; ROM2[3178]<=16'd0; ROM3[3178]<=16'd23806; ROM4[3178]<=16'd57295;
ROM1[3179]<=16'd4817; ROM2[3179]<=16'd0; ROM3[3179]<=16'd23812; ROM4[3179]<=16'd57293;
ROM1[3180]<=16'd4807; ROM2[3180]<=16'd0; ROM3[3180]<=16'd23808; ROM4[3180]<=16'd57287;
ROM1[3181]<=16'd4817; ROM2[3181]<=16'd0; ROM3[3181]<=16'd23797; ROM4[3181]<=16'd57281;
ROM1[3182]<=16'd4846; ROM2[3182]<=16'd0; ROM3[3182]<=16'd23786; ROM4[3182]<=16'd57276;
ROM1[3183]<=16'd4871; ROM2[3183]<=16'd0; ROM3[3183]<=16'd23784; ROM4[3183]<=16'd57282;
ROM1[3184]<=16'd4862; ROM2[3184]<=16'd0; ROM3[3184]<=16'd23791; ROM4[3184]<=16'd57287;
ROM1[3185]<=16'd4834; ROM2[3185]<=16'd0; ROM3[3185]<=16'd23791; ROM4[3185]<=16'd57277;
ROM1[3186]<=16'd4825; ROM2[3186]<=16'd0; ROM3[3186]<=16'd23799; ROM4[3186]<=16'd57280;
ROM1[3187]<=16'd4816; ROM2[3187]<=16'd0; ROM3[3187]<=16'd23806; ROM4[3187]<=16'd57281;
ROM1[3188]<=16'd4818; ROM2[3188]<=16'd0; ROM3[3188]<=16'd23819; ROM4[3188]<=16'd57289;
ROM1[3189]<=16'd4837; ROM2[3189]<=16'd0; ROM3[3189]<=16'd23826; ROM4[3189]<=16'd57303;
ROM1[3190]<=16'd4844; ROM2[3190]<=16'd0; ROM3[3190]<=16'd23800; ROM4[3190]<=16'd57284;
ROM1[3191]<=16'd4855; ROM2[3191]<=16'd0; ROM3[3191]<=16'd23777; ROM4[3191]<=16'd57273;
ROM1[3192]<=16'd4852; ROM2[3192]<=16'd0; ROM3[3192]<=16'd23776; ROM4[3192]<=16'd57275;
ROM1[3193]<=16'd4834; ROM2[3193]<=16'd0; ROM3[3193]<=16'd23780; ROM4[3193]<=16'd57270;
ROM1[3194]<=16'd4836; ROM2[3194]<=16'd0; ROM3[3194]<=16'd23802; ROM4[3194]<=16'd57287;
ROM1[3195]<=16'd4827; ROM2[3195]<=16'd0; ROM3[3195]<=16'd23815; ROM4[3195]<=16'd57293;
ROM1[3196]<=16'd4800; ROM2[3196]<=16'd0; ROM3[3196]<=16'd23803; ROM4[3196]<=16'd57280;
ROM1[3197]<=16'd4797; ROM2[3197]<=16'd0; ROM3[3197]<=16'd23791; ROM4[3197]<=16'd57270;
ROM1[3198]<=16'd4834; ROM2[3198]<=16'd0; ROM3[3198]<=16'd23794; ROM4[3198]<=16'd57274;
ROM1[3199]<=16'd4893; ROM2[3199]<=16'd0; ROM3[3199]<=16'd23803; ROM4[3199]<=16'd57299;
ROM1[3200]<=16'd4888; ROM2[3200]<=16'd0; ROM3[3200]<=16'd23787; ROM4[3200]<=16'd57291;
ROM1[3201]<=16'd4847; ROM2[3201]<=16'd0; ROM3[3201]<=16'd23768; ROM4[3201]<=16'd57271;
ROM1[3202]<=16'd4826; ROM2[3202]<=16'd0; ROM3[3202]<=16'd23780; ROM4[3202]<=16'd57275;
ROM1[3203]<=16'd4817; ROM2[3203]<=16'd0; ROM3[3203]<=16'd23785; ROM4[3203]<=16'd57277;
ROM1[3204]<=16'd4820; ROM2[3204]<=16'd0; ROM3[3204]<=16'd23801; ROM4[3204]<=16'd57290;
ROM1[3205]<=16'd4860; ROM2[3205]<=16'd0; ROM3[3205]<=16'd23839; ROM4[3205]<=16'd57328;
ROM1[3206]<=16'd4880; ROM2[3206]<=16'd0; ROM3[3206]<=16'd23832; ROM4[3206]<=16'd57328;
ROM1[3207]<=16'd4882; ROM2[3207]<=16'd0; ROM3[3207]<=16'd23794; ROM4[3207]<=16'd57301;
ROM1[3208]<=16'd4889; ROM2[3208]<=16'd0; ROM3[3208]<=16'd23780; ROM4[3208]<=16'd57292;
ROM1[3209]<=16'd4865; ROM2[3209]<=16'd0; ROM3[3209]<=16'd23775; ROM4[3209]<=16'd57279;
ROM1[3210]<=16'd4843; ROM2[3210]<=16'd0; ROM3[3210]<=16'd23778; ROM4[3210]<=16'd57275;
ROM1[3211]<=16'd4835; ROM2[3211]<=16'd0; ROM3[3211]<=16'd23791; ROM4[3211]<=16'd57280;
ROM1[3212]<=16'd4830; ROM2[3212]<=16'd0; ROM3[3212]<=16'd23811; ROM4[3212]<=16'd57286;
ROM1[3213]<=16'd4818; ROM2[3213]<=16'd0; ROM3[3213]<=16'd23816; ROM4[3213]<=16'd57283;
ROM1[3214]<=16'd4825; ROM2[3214]<=16'd0; ROM3[3214]<=16'd23811; ROM4[3214]<=16'd57287;
ROM1[3215]<=16'd4873; ROM2[3215]<=16'd0; ROM3[3215]<=16'd23818; ROM4[3215]<=16'd57307;
ROM1[3216]<=16'd4894; ROM2[3216]<=16'd0; ROM3[3216]<=16'd23799; ROM4[3216]<=16'd57300;
ROM1[3217]<=16'd4866; ROM2[3217]<=16'd0; ROM3[3217]<=16'd23773; ROM4[3217]<=16'd57279;
ROM1[3218]<=16'd4848; ROM2[3218]<=16'd0; ROM3[3218]<=16'd23774; ROM4[3218]<=16'd57274;
ROM1[3219]<=16'd4829; ROM2[3219]<=16'd0; ROM3[3219]<=16'd23777; ROM4[3219]<=16'd57269;
ROM1[3220]<=16'd4817; ROM2[3220]<=16'd0; ROM3[3220]<=16'd23787; ROM4[3220]<=16'd57274;
ROM1[3221]<=16'd4813; ROM2[3221]<=16'd0; ROM3[3221]<=16'd23800; ROM4[3221]<=16'd57282;
ROM1[3222]<=16'd4811; ROM2[3222]<=16'd0; ROM3[3222]<=16'd23795; ROM4[3222]<=16'd57278;
ROM1[3223]<=16'd4825; ROM2[3223]<=16'd0; ROM3[3223]<=16'd23780; ROM4[3223]<=16'd57273;
ROM1[3224]<=16'd4852; ROM2[3224]<=16'd0; ROM3[3224]<=16'd23770; ROM4[3224]<=16'd57269;
ROM1[3225]<=16'd4870; ROM2[3225]<=16'd0; ROM3[3225]<=16'd23779; ROM4[3225]<=16'd57283;
ROM1[3226]<=16'd4860; ROM2[3226]<=16'd0; ROM3[3226]<=16'd23789; ROM4[3226]<=16'd57287;
ROM1[3227]<=16'd4842; ROM2[3227]<=16'd0; ROM3[3227]<=16'd23799; ROM4[3227]<=16'd57288;
ROM1[3228]<=16'd4849; ROM2[3228]<=16'd0; ROM3[3228]<=16'd23822; ROM4[3228]<=16'd57309;
ROM1[3229]<=16'd4846; ROM2[3229]<=16'd0; ROM3[3229]<=16'd23839; ROM4[3229]<=16'd57316;
ROM1[3230]<=16'd4821; ROM2[3230]<=16'd0; ROM3[3230]<=16'd23819; ROM4[3230]<=16'd57291;
ROM1[3231]<=16'd4823; ROM2[3231]<=16'd0; ROM3[3231]<=16'd23798; ROM4[3231]<=16'd57275;
ROM1[3232]<=16'd4851; ROM2[3232]<=16'd0; ROM3[3232]<=16'd23782; ROM4[3232]<=16'd57273;
ROM1[3233]<=16'd4865; ROM2[3233]<=16'd0; ROM3[3233]<=16'd23769; ROM4[3233]<=16'd57272;
ROM1[3234]<=16'd4872; ROM2[3234]<=16'd0; ROM3[3234]<=16'd23784; ROM4[3234]<=16'd57290;
ROM1[3235]<=16'd4872; ROM2[3235]<=16'd0; ROM3[3235]<=16'd23802; ROM4[3235]<=16'd57307;
ROM1[3236]<=16'd4859; ROM2[3236]<=16'd0; ROM3[3236]<=16'd23810; ROM4[3236]<=16'd57308;
ROM1[3237]<=16'd4851; ROM2[3237]<=16'd0; ROM3[3237]<=16'd23818; ROM4[3237]<=16'd57314;
ROM1[3238]<=16'd4855; ROM2[3238]<=16'd0; ROM3[3238]<=16'd23832; ROM4[3238]<=16'd57323;
ROM1[3239]<=16'd4842; ROM2[3239]<=16'd0; ROM3[3239]<=16'd23809; ROM4[3239]<=16'd57298;
ROM1[3240]<=16'd4846; ROM2[3240]<=16'd0; ROM3[3240]<=16'd23773; ROM4[3240]<=16'd57273;
ROM1[3241]<=16'd4868; ROM2[3241]<=16'd0; ROM3[3241]<=16'd23759; ROM4[3241]<=16'd57269;
ROM1[3242]<=16'd4861; ROM2[3242]<=16'd0; ROM3[3242]<=16'd23758; ROM4[3242]<=16'd57270;
ROM1[3243]<=16'd4852; ROM2[3243]<=16'd0; ROM3[3243]<=16'd23778; ROM4[3243]<=16'd57286;
ROM1[3244]<=16'd4849; ROM2[3244]<=16'd0; ROM3[3244]<=16'd23798; ROM4[3244]<=16'd57297;
ROM1[3245]<=16'd4833; ROM2[3245]<=16'd0; ROM3[3245]<=16'd23804; ROM4[3245]<=16'd57292;
ROM1[3246]<=16'd4818; ROM2[3246]<=16'd0; ROM3[3246]<=16'd23806; ROM4[3246]<=16'd57291;
ROM1[3247]<=16'd4825; ROM2[3247]<=16'd0; ROM3[3247]<=16'd23810; ROM4[3247]<=16'd57296;
ROM1[3248]<=16'd4850; ROM2[3248]<=16'd0; ROM3[3248]<=16'd23804; ROM4[3248]<=16'd57299;
ROM1[3249]<=16'd4879; ROM2[3249]<=16'd0; ROM3[3249]<=16'd23783; ROM4[3249]<=16'd57294;
ROM1[3250]<=16'd4886; ROM2[3250]<=16'd0; ROM3[3250]<=16'd23782; ROM4[3250]<=16'd57297;
ROM1[3251]<=16'd4880; ROM2[3251]<=16'd0; ROM3[3251]<=16'd23796; ROM4[3251]<=16'd57309;
ROM1[3252]<=16'd4856; ROM2[3252]<=16'd0; ROM3[3252]<=16'd23803; ROM4[3252]<=16'd57307;
ROM1[3253]<=16'd4845; ROM2[3253]<=16'd0; ROM3[3253]<=16'd23812; ROM4[3253]<=16'd57313;
ROM1[3254]<=16'd4818; ROM2[3254]<=16'd0; ROM3[3254]<=16'd23804; ROM4[3254]<=16'd57303;
ROM1[3255]<=16'd4804; ROM2[3255]<=16'd0; ROM3[3255]<=16'd23789; ROM4[3255]<=16'd57286;
ROM1[3256]<=16'd4833; ROM2[3256]<=16'd0; ROM3[3256]<=16'd23787; ROM4[3256]<=16'd57291;
ROM1[3257]<=16'd4857; ROM2[3257]<=16'd0; ROM3[3257]<=16'd23771; ROM4[3257]<=16'd57284;
ROM1[3258]<=16'd4881; ROM2[3258]<=16'd0; ROM3[3258]<=16'd23767; ROM4[3258]<=16'd57289;
ROM1[3259]<=16'd4870; ROM2[3259]<=16'd0; ROM3[3259]<=16'd23766; ROM4[3259]<=16'd57284;
ROM1[3260]<=16'd4839; ROM2[3260]<=16'd0; ROM3[3260]<=16'd23761; ROM4[3260]<=16'd57270;
ROM1[3261]<=16'd4837; ROM2[3261]<=16'd0; ROM3[3261]<=16'd23783; ROM4[3261]<=16'd57287;
ROM1[3262]<=16'd4817; ROM2[3262]<=16'd0; ROM3[3262]<=16'd23786; ROM4[3262]<=16'd57287;
ROM1[3263]<=16'd4791; ROM2[3263]<=16'd0; ROM3[3263]<=16'd23769; ROM4[3263]<=16'd57265;
ROM1[3264]<=16'd4811; ROM2[3264]<=16'd0; ROM3[3264]<=16'd23771; ROM4[3264]<=16'd57272;
ROM1[3265]<=16'd4843; ROM2[3265]<=16'd0; ROM3[3265]<=16'd23761; ROM4[3265]<=16'd57272;
ROM1[3266]<=16'd4871; ROM2[3266]<=16'd0; ROM3[3266]<=16'd23757; ROM4[3266]<=16'd57274;
ROM1[3267]<=16'd4879; ROM2[3267]<=16'd0; ROM3[3267]<=16'd23773; ROM4[3267]<=16'd57293;
ROM1[3268]<=16'd4861; ROM2[3268]<=16'd0; ROM3[3268]<=16'd23778; ROM4[3268]<=16'd57295;
ROM1[3269]<=16'd4838; ROM2[3269]<=16'd0; ROM3[3269]<=16'd23777; ROM4[3269]<=16'd57289;
ROM1[3270]<=16'd4827; ROM2[3270]<=16'd0; ROM3[3270]<=16'd23783; ROM4[3270]<=16'd57293;
ROM1[3271]<=16'd4824; ROM2[3271]<=16'd0; ROM3[3271]<=16'd23799; ROM4[3271]<=16'd57300;
ROM1[3272]<=16'd4834; ROM2[3272]<=16'd0; ROM3[3272]<=16'd23807; ROM4[3272]<=16'd57310;
ROM1[3273]<=16'd4861; ROM2[3273]<=16'd0; ROM3[3273]<=16'd23800; ROM4[3273]<=16'd57315;
ROM1[3274]<=16'd4895; ROM2[3274]<=16'd0; ROM3[3274]<=16'd23790; ROM4[3274]<=16'd57314;
ROM1[3275]<=16'd4899; ROM2[3275]<=16'd0; ROM3[3275]<=16'd23787; ROM4[3275]<=16'd57315;
ROM1[3276]<=16'd4888; ROM2[3276]<=16'd0; ROM3[3276]<=16'd23796; ROM4[3276]<=16'd57322;
ROM1[3277]<=16'd4881; ROM2[3277]<=16'd0; ROM3[3277]<=16'd23817; ROM4[3277]<=16'd57334;
ROM1[3278]<=16'd4865; ROM2[3278]<=16'd0; ROM3[3278]<=16'd23826; ROM4[3278]<=16'd57334;
ROM1[3279]<=16'd4844; ROM2[3279]<=16'd0; ROM3[3279]<=16'd23822; ROM4[3279]<=16'd57324;
ROM1[3280]<=16'd4839; ROM2[3280]<=16'd0; ROM3[3280]<=16'd23818; ROM4[3280]<=16'd57317;
ROM1[3281]<=16'd4844; ROM2[3281]<=16'd0; ROM3[3281]<=16'd23803; ROM4[3281]<=16'd57306;
ROM1[3282]<=16'd4871; ROM2[3282]<=16'd0; ROM3[3282]<=16'd23790; ROM4[3282]<=16'd57301;
ROM1[3283]<=16'd4894; ROM2[3283]<=16'd0; ROM3[3283]<=16'd23790; ROM4[3283]<=16'd57309;
ROM1[3284]<=16'd4883; ROM2[3284]<=16'd0; ROM3[3284]<=16'd23795; ROM4[3284]<=16'd57315;
ROM1[3285]<=16'd4871; ROM2[3285]<=16'd0; ROM3[3285]<=16'd23808; ROM4[3285]<=16'd57323;
ROM1[3286]<=16'd4866; ROM2[3286]<=16'd0; ROM3[3286]<=16'd23823; ROM4[3286]<=16'd57331;
ROM1[3287]<=16'd4852; ROM2[3287]<=16'd0; ROM3[3287]<=16'd23833; ROM4[3287]<=16'd57331;
ROM1[3288]<=16'd4832; ROM2[3288]<=16'd0; ROM3[3288]<=16'd23832; ROM4[3288]<=16'd57324;
ROM1[3289]<=16'd4831; ROM2[3289]<=16'd0; ROM3[3289]<=16'd23823; ROM4[3289]<=16'd57314;
ROM1[3290]<=16'd4863; ROM2[3290]<=16'd0; ROM3[3290]<=16'd23813; ROM4[3290]<=16'd57313;
ROM1[3291]<=16'd4894; ROM2[3291]<=16'd0; ROM3[3291]<=16'd23809; ROM4[3291]<=16'd57324;
ROM1[3292]<=16'd4886; ROM2[3292]<=16'd0; ROM3[3292]<=16'd23813; ROM4[3292]<=16'd57321;
ROM1[3293]<=16'd4868; ROM2[3293]<=16'd0; ROM3[3293]<=16'd23812; ROM4[3293]<=16'd57315;
ROM1[3294]<=16'd4852; ROM2[3294]<=16'd0; ROM3[3294]<=16'd23816; ROM4[3294]<=16'd57312;
ROM1[3295]<=16'd4849; ROM2[3295]<=16'd0; ROM3[3295]<=16'd23834; ROM4[3295]<=16'd57319;
ROM1[3296]<=16'd4843; ROM2[3296]<=16'd0; ROM3[3296]<=16'd23833; ROM4[3296]<=16'd57317;
ROM1[3297]<=16'd4832; ROM2[3297]<=16'd0; ROM3[3297]<=16'd23810; ROM4[3297]<=16'd57299;
ROM1[3298]<=16'd4859; ROM2[3298]<=16'd0; ROM3[3298]<=16'd23806; ROM4[3298]<=16'd57307;
ROM1[3299]<=16'd4892; ROM2[3299]<=16'd0; ROM3[3299]<=16'd23793; ROM4[3299]<=16'd57310;
ROM1[3300]<=16'd4895; ROM2[3300]<=16'd0; ROM3[3300]<=16'd23788; ROM4[3300]<=16'd57307;
ROM1[3301]<=16'd4881; ROM2[3301]<=16'd0; ROM3[3301]<=16'd23797; ROM4[3301]<=16'd57311;
ROM1[3302]<=16'd4859; ROM2[3302]<=16'd0; ROM3[3302]<=16'd23800; ROM4[3302]<=16'd57304;
ROM1[3303]<=16'd4842; ROM2[3303]<=16'd0; ROM3[3303]<=16'd23797; ROM4[3303]<=16'd57296;
ROM1[3304]<=16'd4833; ROM2[3304]<=16'd0; ROM3[3304]<=16'd23803; ROM4[3304]<=16'd57296;
ROM1[3305]<=16'd4844; ROM2[3305]<=16'd0; ROM3[3305]<=16'd23818; ROM4[3305]<=16'd57307;
ROM1[3306]<=16'd4865; ROM2[3306]<=16'd0; ROM3[3306]<=16'd23818; ROM4[3306]<=16'd57310;
ROM1[3307]<=16'd4898; ROM2[3307]<=16'd0; ROM3[3307]<=16'd23804; ROM4[3307]<=16'd57307;
ROM1[3308]<=16'd4906; ROM2[3308]<=16'd0; ROM3[3308]<=16'd23793; ROM4[3308]<=16'd57303;
ROM1[3309]<=16'd4891; ROM2[3309]<=16'd0; ROM3[3309]<=16'd23797; ROM4[3309]<=16'd57302;
ROM1[3310]<=16'd4882; ROM2[3310]<=16'd0; ROM3[3310]<=16'd23813; ROM4[3310]<=16'd57311;
ROM1[3311]<=16'd4863; ROM2[3311]<=16'd0; ROM3[3311]<=16'd23820; ROM4[3311]<=16'd57311;
ROM1[3312]<=16'd4844; ROM2[3312]<=16'd0; ROM3[3312]<=16'd23819; ROM4[3312]<=16'd57304;
ROM1[3313]<=16'd4840; ROM2[3313]<=16'd0; ROM3[3313]<=16'd23825; ROM4[3313]<=16'd57304;
ROM1[3314]<=16'd4850; ROM2[3314]<=16'd0; ROM3[3314]<=16'd23823; ROM4[3314]<=16'd57303;
ROM1[3315]<=16'd4874; ROM2[3315]<=16'd0; ROM3[3315]<=16'd23812; ROM4[3315]<=16'd57302;
ROM1[3316]<=16'd4892; ROM2[3316]<=16'd0; ROM3[3316]<=16'd23801; ROM4[3316]<=16'd57302;
ROM1[3317]<=16'd4885; ROM2[3317]<=16'd0; ROM3[3317]<=16'd23801; ROM4[3317]<=16'd57300;
ROM1[3318]<=16'd4860; ROM2[3318]<=16'd0; ROM3[3318]<=16'd23803; ROM4[3318]<=16'd57291;
ROM1[3319]<=16'd4847; ROM2[3319]<=16'd0; ROM3[3319]<=16'd23809; ROM4[3319]<=16'd57285;
ROM1[3320]<=16'd4851; ROM2[3320]<=16'd0; ROM3[3320]<=16'd23826; ROM4[3320]<=16'd57298;
ROM1[3321]<=16'd4853; ROM2[3321]<=16'd0; ROM3[3321]<=16'd23839; ROM4[3321]<=16'd57310;
ROM1[3322]<=16'd4863; ROM2[3322]<=16'd0; ROM3[3322]<=16'd23841; ROM4[3322]<=16'd57319;
ROM1[3323]<=16'd4869; ROM2[3323]<=16'd0; ROM3[3323]<=16'd23816; ROM4[3323]<=16'd57305;
ROM1[3324]<=16'd4892; ROM2[3324]<=16'd0; ROM3[3324]<=16'd23793; ROM4[3324]<=16'd57293;
ROM1[3325]<=16'd4907; ROM2[3325]<=16'd0; ROM3[3325]<=16'd23793; ROM4[3325]<=16'd57302;
ROM1[3326]<=16'd4877; ROM2[3326]<=16'd0; ROM3[3326]<=16'd23782; ROM4[3326]<=16'd57285;
ROM1[3327]<=16'd4856; ROM2[3327]<=16'd0; ROM3[3327]<=16'd23791; ROM4[3327]<=16'd57286;
ROM1[3328]<=16'd4848; ROM2[3328]<=16'd0; ROM3[3328]<=16'd23806; ROM4[3328]<=16'd57295;
ROM1[3329]<=16'd4821; ROM2[3329]<=16'd0; ROM3[3329]<=16'd23803; ROM4[3329]<=16'd57284;
ROM1[3330]<=16'd4820; ROM2[3330]<=16'd0; ROM3[3330]<=16'd23807; ROM4[3330]<=16'd57286;
ROM1[3331]<=16'd4858; ROM2[3331]<=16'd0; ROM3[3331]<=16'd23817; ROM4[3331]<=16'd57304;
ROM1[3332]<=16'd4894; ROM2[3332]<=16'd0; ROM3[3332]<=16'd23807; ROM4[3332]<=16'd57306;
ROM1[3333]<=16'd4886; ROM2[3333]<=16'd0; ROM3[3333]<=16'd23776; ROM4[3333]<=16'd57283;
ROM1[3334]<=16'd4863; ROM2[3334]<=16'd0; ROM3[3334]<=16'd23769; ROM4[3334]<=16'd57275;
ROM1[3335]<=16'd4850; ROM2[3335]<=16'd0; ROM3[3335]<=16'd23786; ROM4[3335]<=16'd57283;
ROM1[3336]<=16'd4840; ROM2[3336]<=16'd0; ROM3[3336]<=16'd23799; ROM4[3336]<=16'd57287;
ROM1[3337]<=16'd4828; ROM2[3337]<=16'd0; ROM3[3337]<=16'd23807; ROM4[3337]<=16'd57284;
ROM1[3338]<=16'd4825; ROM2[3338]<=16'd0; ROM3[3338]<=16'd23813; ROM4[3338]<=16'd57287;
ROM1[3339]<=16'd4836; ROM2[3339]<=16'd0; ROM3[3339]<=16'd23806; ROM4[3339]<=16'd57286;
ROM1[3340]<=16'd4866; ROM2[3340]<=16'd0; ROM3[3340]<=16'd23799; ROM4[3340]<=16'd57290;
ROM1[3341]<=16'd4901; ROM2[3341]<=16'd0; ROM3[3341]<=16'd23800; ROM4[3341]<=16'd57304;
ROM1[3342]<=16'd4902; ROM2[3342]<=16'd0; ROM3[3342]<=16'd23803; ROM4[3342]<=16'd57309;
ROM1[3343]<=16'd4885; ROM2[3343]<=16'd0; ROM3[3343]<=16'd23807; ROM4[3343]<=16'd57309;
ROM1[3344]<=16'd4880; ROM2[3344]<=16'd0; ROM3[3344]<=16'd23822; ROM4[3344]<=16'd57317;
ROM1[3345]<=16'd4874; ROM2[3345]<=16'd0; ROM3[3345]<=16'd23839; ROM4[3345]<=16'd57331;
ROM1[3346]<=16'd4859; ROM2[3346]<=16'd0; ROM3[3346]<=16'd23849; ROM4[3346]<=16'd57334;
ROM1[3347]<=16'd4868; ROM2[3347]<=16'd0; ROM3[3347]<=16'd23854; ROM4[3347]<=16'd57337;
ROM1[3348]<=16'd4887; ROM2[3348]<=16'd0; ROM3[3348]<=16'd23842; ROM4[3348]<=16'd57337;
ROM1[3349]<=16'd4913; ROM2[3349]<=16'd0; ROM3[3349]<=16'd23825; ROM4[3349]<=16'd57333;
ROM1[3350]<=16'd4912; ROM2[3350]<=16'd0; ROM3[3350]<=16'd23814; ROM4[3350]<=16'd57326;
ROM1[3351]<=16'd4881; ROM2[3351]<=16'd0; ROM3[3351]<=16'd23811; ROM4[3351]<=16'd57320;
ROM1[3352]<=16'd4857; ROM2[3352]<=16'd0; ROM3[3352]<=16'd23822; ROM4[3352]<=16'd57321;
ROM1[3353]<=16'd4850; ROM2[3353]<=16'd0; ROM3[3353]<=16'd23836; ROM4[3353]<=16'd57326;
ROM1[3354]<=16'd4841; ROM2[3354]<=16'd0; ROM3[3354]<=16'd23846; ROM4[3354]<=16'd57330;
ROM1[3355]<=16'd4844; ROM2[3355]<=16'd0; ROM3[3355]<=16'd23852; ROM4[3355]<=16'd57333;
ROM1[3356]<=16'd4865; ROM2[3356]<=16'd0; ROM3[3356]<=16'd23848; ROM4[3356]<=16'd57338;
ROM1[3357]<=16'd4895; ROM2[3357]<=16'd0; ROM3[3357]<=16'd23841; ROM4[3357]<=16'd57342;
ROM1[3358]<=16'd4902; ROM2[3358]<=16'd0; ROM3[3358]<=16'd23827; ROM4[3358]<=16'd57338;
ROM1[3359]<=16'd4884; ROM2[3359]<=16'd0; ROM3[3359]<=16'd23828; ROM4[3359]<=16'd57333;
ROM1[3360]<=16'd4870; ROM2[3360]<=16'd0; ROM3[3360]<=16'd23838; ROM4[3360]<=16'd57334;
ROM1[3361]<=16'd4848; ROM2[3361]<=16'd0; ROM3[3361]<=16'd23836; ROM4[3361]<=16'd57328;
ROM1[3362]<=16'd4819; ROM2[3362]<=16'd0; ROM3[3362]<=16'd23835; ROM4[3362]<=16'd57317;
ROM1[3363]<=16'd4816; ROM2[3363]<=16'd0; ROM3[3363]<=16'd23842; ROM4[3363]<=16'd57319;
ROM1[3364]<=16'd4817; ROM2[3364]<=16'd0; ROM3[3364]<=16'd23828; ROM4[3364]<=16'd57314;
ROM1[3365]<=16'd4843; ROM2[3365]<=16'd0; ROM3[3365]<=16'd23811; ROM4[3365]<=16'd57310;
ROM1[3366]<=16'd4884; ROM2[3366]<=16'd0; ROM3[3366]<=16'd23808; ROM4[3366]<=16'd57319;
ROM1[3367]<=16'd4877; ROM2[3367]<=16'd0; ROM3[3367]<=16'd23806; ROM4[3367]<=16'd57317;
ROM1[3368]<=16'd4849; ROM2[3368]<=16'd0; ROM3[3368]<=16'd23806; ROM4[3368]<=16'd57309;
ROM1[3369]<=16'd4837; ROM2[3369]<=16'd0; ROM3[3369]<=16'd23820; ROM4[3369]<=16'd57313;
ROM1[3370]<=16'd4839; ROM2[3370]<=16'd0; ROM3[3370]<=16'd23840; ROM4[3370]<=16'd57330;
ROM1[3371]<=16'd4822; ROM2[3371]<=16'd0; ROM3[3371]<=16'd23835; ROM4[3371]<=16'd57324;
ROM1[3372]<=16'd4822; ROM2[3372]<=16'd0; ROM3[3372]<=16'd23827; ROM4[3372]<=16'd57315;
ROM1[3373]<=16'd4850; ROM2[3373]<=16'd0; ROM3[3373]<=16'd23821; ROM4[3373]<=16'd57319;
ROM1[3374]<=16'd4891; ROM2[3374]<=16'd0; ROM3[3374]<=16'd23813; ROM4[3374]<=16'd57322;
ROM1[3375]<=16'd4885; ROM2[3375]<=16'd0; ROM3[3375]<=16'd23808; ROM4[3375]<=16'd57319;
ROM1[3376]<=16'd4869; ROM2[3376]<=16'd0; ROM3[3376]<=16'd23811; ROM4[3376]<=16'd57318;
ROM1[3377]<=16'd4856; ROM2[3377]<=16'd0; ROM3[3377]<=16'd23816; ROM4[3377]<=16'd57314;
ROM1[3378]<=16'd4830; ROM2[3378]<=16'd0; ROM3[3378]<=16'd23814; ROM4[3378]<=16'd57305;
ROM1[3379]<=16'd4819; ROM2[3379]<=16'd0; ROM3[3379]<=16'd23818; ROM4[3379]<=16'd57303;
ROM1[3380]<=16'd4819; ROM2[3380]<=16'd0; ROM3[3380]<=16'd23823; ROM4[3380]<=16'd57308;
ROM1[3381]<=16'd4839; ROM2[3381]<=16'd0; ROM3[3381]<=16'd23825; ROM4[3381]<=16'd57322;
ROM1[3382]<=16'd4873; ROM2[3382]<=16'd0; ROM3[3382]<=16'd23810; ROM4[3382]<=16'd57320;
ROM1[3383]<=16'd4892; ROM2[3383]<=16'd0; ROM3[3383]<=16'd23804; ROM4[3383]<=16'd57319;
ROM1[3384]<=16'd4885; ROM2[3384]<=16'd0; ROM3[3384]<=16'd23810; ROM4[3384]<=16'd57325;
ROM1[3385]<=16'd4865; ROM2[3385]<=16'd0; ROM3[3385]<=16'd23812; ROM4[3385]<=16'd57323;
ROM1[3386]<=16'd4848; ROM2[3386]<=16'd0; ROM3[3386]<=16'd23820; ROM4[3386]<=16'd57322;
ROM1[3387]<=16'd4834; ROM2[3387]<=16'd0; ROM3[3387]<=16'd23830; ROM4[3387]<=16'd57329;
ROM1[3388]<=16'd4819; ROM2[3388]<=16'd0; ROM3[3388]<=16'd23829; ROM4[3388]<=16'd57324;
ROM1[3389]<=16'd4822; ROM2[3389]<=16'd0; ROM3[3389]<=16'd23819; ROM4[3389]<=16'd57313;
ROM1[3390]<=16'd4849; ROM2[3390]<=16'd0; ROM3[3390]<=16'd23806; ROM4[3390]<=16'd57312;
ROM1[3391]<=16'd4880; ROM2[3391]<=16'd0; ROM3[3391]<=16'd23794; ROM4[3391]<=16'd57315;
ROM1[3392]<=16'd4883; ROM2[3392]<=16'd0; ROM3[3392]<=16'd23797; ROM4[3392]<=16'd57318;
ROM1[3393]<=16'd4871; ROM2[3393]<=16'd0; ROM3[3393]<=16'd23811; ROM4[3393]<=16'd57321;
ROM1[3394]<=16'd4855; ROM2[3394]<=16'd0; ROM3[3394]<=16'd23821; ROM4[3394]<=16'd57323;
ROM1[3395]<=16'd4846; ROM2[3395]<=16'd0; ROM3[3395]<=16'd23836; ROM4[3395]<=16'd57332;
ROM1[3396]<=16'd4849; ROM2[3396]<=16'd0; ROM3[3396]<=16'd23853; ROM4[3396]<=16'd57340;
ROM1[3397]<=16'd4864; ROM2[3397]<=16'd0; ROM3[3397]<=16'd23860; ROM4[3397]<=16'd57349;
ROM1[3398]<=16'd4897; ROM2[3398]<=16'd0; ROM3[3398]<=16'd23863; ROM4[3398]<=16'd57358;
ROM1[3399]<=16'd4908; ROM2[3399]<=16'd0; ROM3[3399]<=16'd23834; ROM4[3399]<=16'd57341;
ROM1[3400]<=16'd4898; ROM2[3400]<=16'd0; ROM3[3400]<=16'd23816; ROM4[3400]<=16'd57327;
ROM1[3401]<=16'd4886; ROM2[3401]<=16'd0; ROM3[3401]<=16'd23828; ROM4[3401]<=16'd57335;
ROM1[3402]<=16'd4865; ROM2[3402]<=16'd0; ROM3[3402]<=16'd23835; ROM4[3402]<=16'd57335;
ROM1[3403]<=16'd4857; ROM2[3403]<=16'd0; ROM3[3403]<=16'd23844; ROM4[3403]<=16'd57335;
ROM1[3404]<=16'd4848; ROM2[3404]<=16'd0; ROM3[3404]<=16'd23857; ROM4[3404]<=16'd57345;
ROM1[3405]<=16'd4840; ROM2[3405]<=16'd0; ROM3[3405]<=16'd23848; ROM4[3405]<=16'd57337;
ROM1[3406]<=16'd4850; ROM2[3406]<=16'd0; ROM3[3406]<=16'd23834; ROM4[3406]<=16'd57325;
ROM1[3407]<=16'd4887; ROM2[3407]<=16'd0; ROM3[3407]<=16'd23826; ROM4[3407]<=16'd57330;
ROM1[3408]<=16'd4898; ROM2[3408]<=16'd0; ROM3[3408]<=16'd23816; ROM4[3408]<=16'd57328;
ROM1[3409]<=16'd4878; ROM2[3409]<=16'd0; ROM3[3409]<=16'd23815; ROM4[3409]<=16'd57322;
ROM1[3410]<=16'd4866; ROM2[3410]<=16'd0; ROM3[3410]<=16'd23825; ROM4[3410]<=16'd57327;
ROM1[3411]<=16'd4856; ROM2[3411]<=16'd0; ROM3[3411]<=16'd23838; ROM4[3411]<=16'd57333;
ROM1[3412]<=16'd4839; ROM2[3412]<=16'd0; ROM3[3412]<=16'd23842; ROM4[3412]<=16'd57332;
ROM1[3413]<=16'd4830; ROM2[3413]<=16'd0; ROM3[3413]<=16'd23844; ROM4[3413]<=16'd57327;
ROM1[3414]<=16'd4847; ROM2[3414]<=16'd0; ROM3[3414]<=16'd23846; ROM4[3414]<=16'd57335;
ROM1[3415]<=16'd4900; ROM2[3415]<=16'd0; ROM3[3415]<=16'd23862; ROM4[3415]<=16'd57366;
ROM1[3416]<=16'd4936; ROM2[3416]<=16'd0; ROM3[3416]<=16'd23863; ROM4[3416]<=16'd57374;
ROM1[3417]<=16'd4908; ROM2[3417]<=16'd0; ROM3[3417]<=16'd23842; ROM4[3417]<=16'd57355;
ROM1[3418]<=16'd4887; ROM2[3418]<=16'd0; ROM3[3418]<=16'd23851; ROM4[3418]<=16'd57356;
ROM1[3419]<=16'd4878; ROM2[3419]<=16'd0; ROM3[3419]<=16'd23870; ROM4[3419]<=16'd57362;
ROM1[3420]<=16'd4856; ROM2[3420]<=16'd0; ROM3[3420]<=16'd23867; ROM4[3420]<=16'd57356;
ROM1[3421]<=16'd4841; ROM2[3421]<=16'd0; ROM3[3421]<=16'd23868; ROM4[3421]<=16'd57348;
ROM1[3422]<=16'd4840; ROM2[3422]<=16'd0; ROM3[3422]<=16'd23861; ROM4[3422]<=16'd57341;
ROM1[3423]<=16'd4862; ROM2[3423]<=16'd0; ROM3[3423]<=16'd23847; ROM4[3423]<=16'd57337;
ROM1[3424]<=16'd4895; ROM2[3424]<=16'd0; ROM3[3424]<=16'd23838; ROM4[3424]<=16'd57339;
ROM1[3425]<=16'd4910; ROM2[3425]<=16'd0; ROM3[3425]<=16'd23843; ROM4[3425]<=16'd57349;
ROM1[3426]<=16'd4902; ROM2[3426]<=16'd0; ROM3[3426]<=16'd23855; ROM4[3426]<=16'd57356;
ROM1[3427]<=16'd4880; ROM2[3427]<=16'd0; ROM3[3427]<=16'd23859; ROM4[3427]<=16'd57353;
ROM1[3428]<=16'd4872; ROM2[3428]<=16'd0; ROM3[3428]<=16'd23871; ROM4[3428]<=16'd57362;
ROM1[3429]<=16'd4864; ROM2[3429]<=16'd0; ROM3[3429]<=16'd23883; ROM4[3429]<=16'd57367;
ROM1[3430]<=16'd4864; ROM2[3430]<=16'd0; ROM3[3430]<=16'd23879; ROM4[3430]<=16'd57362;
ROM1[3431]<=16'd4871; ROM2[3431]<=16'd0; ROM3[3431]<=16'd23863; ROM4[3431]<=16'd57353;
ROM1[3432]<=16'd4894; ROM2[3432]<=16'd0; ROM3[3432]<=16'd23845; ROM4[3432]<=16'd57345;
ROM1[3433]<=16'd4910; ROM2[3433]<=16'd0; ROM3[3433]<=16'd23843; ROM4[3433]<=16'd57351;
ROM1[3434]<=16'd4898; ROM2[3434]<=16'd0; ROM3[3434]<=16'd23848; ROM4[3434]<=16'd57354;
ROM1[3435]<=16'd4875; ROM2[3435]<=16'd0; ROM3[3435]<=16'd23850; ROM4[3435]<=16'd57347;
ROM1[3436]<=16'd4862; ROM2[3436]<=16'd0; ROM3[3436]<=16'd23858; ROM4[3436]<=16'd57349;
ROM1[3437]<=16'd4861; ROM2[3437]<=16'd0; ROM3[3437]<=16'd23880; ROM4[3437]<=16'd57362;
ROM1[3438]<=16'd4850; ROM2[3438]<=16'd0; ROM3[3438]<=16'd23881; ROM4[3438]<=16'd57363;
ROM1[3439]<=16'd4863; ROM2[3439]<=16'd0; ROM3[3439]<=16'd23878; ROM4[3439]<=16'd57363;
ROM1[3440]<=16'd4907; ROM2[3440]<=16'd0; ROM3[3440]<=16'd23877; ROM4[3440]<=16'd57374;
ROM1[3441]<=16'd4915; ROM2[3441]<=16'd0; ROM3[3441]<=16'd23846; ROM4[3441]<=16'd57355;
ROM1[3442]<=16'd4903; ROM2[3442]<=16'd0; ROM3[3442]<=16'd23838; ROM4[3442]<=16'd57346;
ROM1[3443]<=16'd4895; ROM2[3443]<=16'd0; ROM3[3443]<=16'd23851; ROM4[3443]<=16'd57353;
ROM1[3444]<=16'd4866; ROM2[3444]<=16'd0; ROM3[3444]<=16'd23847; ROM4[3444]<=16'd57341;
ROM1[3445]<=16'd4845; ROM2[3445]<=16'd0; ROM3[3445]<=16'd23850; ROM4[3445]<=16'd57339;
ROM1[3446]<=16'd4837; ROM2[3446]<=16'd0; ROM3[3446]<=16'd23859; ROM4[3446]<=16'd57345;
ROM1[3447]<=16'd4835; ROM2[3447]<=16'd0; ROM3[3447]<=16'd23854; ROM4[3447]<=16'd57343;
ROM1[3448]<=16'd4858; ROM2[3448]<=16'd0; ROM3[3448]<=16'd23841; ROM4[3448]<=16'd57338;
ROM1[3449]<=16'd4900; ROM2[3449]<=16'd0; ROM3[3449]<=16'd23838; ROM4[3449]<=16'd57344;
ROM1[3450]<=16'd4912; ROM2[3450]<=16'd0; ROM3[3450]<=16'd23851; ROM4[3450]<=16'd57351;
ROM1[3451]<=16'd4888; ROM2[3451]<=16'd0; ROM3[3451]<=16'd23850; ROM4[3451]<=16'd57346;
ROM1[3452]<=16'd4869; ROM2[3452]<=16'd0; ROM3[3452]<=16'd23858; ROM4[3452]<=16'd57348;
ROM1[3453]<=16'd4860; ROM2[3453]<=16'd0; ROM3[3453]<=16'd23868; ROM4[3453]<=16'd57353;
ROM1[3454]<=16'd4847; ROM2[3454]<=16'd0; ROM3[3454]<=16'd23869; ROM4[3454]<=16'd57353;
ROM1[3455]<=16'd4844; ROM2[3455]<=16'd0; ROM3[3455]<=16'd23869; ROM4[3455]<=16'd57346;
ROM1[3456]<=16'd4850; ROM2[3456]<=16'd0; ROM3[3456]<=16'd23853; ROM4[3456]<=16'd57333;
ROM1[3457]<=16'd4883; ROM2[3457]<=16'd0; ROM3[3457]<=16'd23842; ROM4[3457]<=16'd57335;
ROM1[3458]<=16'd4894; ROM2[3458]<=16'd0; ROM3[3458]<=16'd23833; ROM4[3458]<=16'd57331;
ROM1[3459]<=16'd4881; ROM2[3459]<=16'd0; ROM3[3459]<=16'd23833; ROM4[3459]<=16'd57330;
ROM1[3460]<=16'd4861; ROM2[3460]<=16'd0; ROM3[3460]<=16'd23842; ROM4[3460]<=16'd57330;
ROM1[3461]<=16'd4846; ROM2[3461]<=16'd0; ROM3[3461]<=16'd23845; ROM4[3461]<=16'd57328;
ROM1[3462]<=16'd4837; ROM2[3462]<=16'd0; ROM3[3462]<=16'd23850; ROM4[3462]<=16'd57332;
ROM1[3463]<=16'd4841; ROM2[3463]<=16'd0; ROM3[3463]<=16'd23863; ROM4[3463]<=16'd57342;
ROM1[3464]<=16'd4868; ROM2[3464]<=16'd0; ROM3[3464]<=16'd23871; ROM4[3464]<=16'd57353;
ROM1[3465]<=16'd4895; ROM2[3465]<=16'd0; ROM3[3465]<=16'd23861; ROM4[3465]<=16'd57350;
ROM1[3466]<=16'd4910; ROM2[3466]<=16'd0; ROM3[3466]<=16'd23847; ROM4[3466]<=16'd57343;
ROM1[3467]<=16'd4905; ROM2[3467]<=16'd0; ROM3[3467]<=16'd23850; ROM4[3467]<=16'd57349;
ROM1[3468]<=16'd4889; ROM2[3468]<=16'd0; ROM3[3468]<=16'd23857; ROM4[3468]<=16'd57352;
ROM1[3469]<=16'd4861; ROM2[3469]<=16'd0; ROM3[3469]<=16'd23848; ROM4[3469]<=16'd57338;
ROM1[3470]<=16'd4849; ROM2[3470]<=16'd0; ROM3[3470]<=16'd23841; ROM4[3470]<=16'd57332;
ROM1[3471]<=16'd4839; ROM2[3471]<=16'd0; ROM3[3471]<=16'd23845; ROM4[3471]<=16'd57330;
ROM1[3472]<=16'd4843; ROM2[3472]<=16'd0; ROM3[3472]<=16'd23843; ROM4[3472]<=16'd57328;
ROM1[3473]<=16'd4868; ROM2[3473]<=16'd0; ROM3[3473]<=16'd23835; ROM4[3473]<=16'd57329;
ROM1[3474]<=16'd4889; ROM2[3474]<=16'd0; ROM3[3474]<=16'd23820; ROM4[3474]<=16'd57322;
ROM1[3475]<=16'd4897; ROM2[3475]<=16'd0; ROM3[3475]<=16'd23820; ROM4[3475]<=16'd57327;
ROM1[3476]<=16'd4880; ROM2[3476]<=16'd0; ROM3[3476]<=16'd23828; ROM4[3476]<=16'd57325;
ROM1[3477]<=16'd4849; ROM2[3477]<=16'd0; ROM3[3477]<=16'd23829; ROM4[3477]<=16'd57317;
ROM1[3478]<=16'd4837; ROM2[3478]<=16'd0; ROM3[3478]<=16'd23835; ROM4[3478]<=16'd57321;
ROM1[3479]<=16'd4824; ROM2[3479]<=16'd0; ROM3[3479]<=16'd23839; ROM4[3479]<=16'd57319;
ROM1[3480]<=16'd4815; ROM2[3480]<=16'd0; ROM3[3480]<=16'd23834; ROM4[3480]<=16'd57312;
ROM1[3481]<=16'd4839; ROM2[3481]<=16'd0; ROM3[3481]<=16'd23836; ROM4[3481]<=16'd57318;
ROM1[3482]<=16'd4873; ROM2[3482]<=16'd0; ROM3[3482]<=16'd23828; ROM4[3482]<=16'd57323;
ROM1[3483]<=16'd4896; ROM2[3483]<=16'd0; ROM3[3483]<=16'd23832; ROM4[3483]<=16'd57338;
ROM1[3484]<=16'd4891; ROM2[3484]<=16'd0; ROM3[3484]<=16'd23844; ROM4[3484]<=16'd57348;
ROM1[3485]<=16'd4884; ROM2[3485]<=16'd0; ROM3[3485]<=16'd23860; ROM4[3485]<=16'd57358;
ROM1[3486]<=16'd4875; ROM2[3486]<=16'd0; ROM3[3486]<=16'd23876; ROM4[3486]<=16'd57364;
ROM1[3487]<=16'd4833; ROM2[3487]<=16'd0; ROM3[3487]<=16'd23853; ROM4[3487]<=16'd57334;
ROM1[3488]<=16'd4828; ROM2[3488]<=16'd0; ROM3[3488]<=16'd23849; ROM4[3488]<=16'd57331;
ROM1[3489]<=16'd4846; ROM2[3489]<=16'd0; ROM3[3489]<=16'd23851; ROM4[3489]<=16'd57336;
ROM1[3490]<=16'd4862; ROM2[3490]<=16'd0; ROM3[3490]<=16'd23831; ROM4[3490]<=16'd57326;
ROM1[3491]<=16'd4886; ROM2[3491]<=16'd0; ROM3[3491]<=16'd23818; ROM4[3491]<=16'd57323;
ROM1[3492]<=16'd4880; ROM2[3492]<=16'd0; ROM3[3492]<=16'd23816; ROM4[3492]<=16'd57323;
ROM1[3493]<=16'd4870; ROM2[3493]<=16'd0; ROM3[3493]<=16'd23829; ROM4[3493]<=16'd57328;
ROM1[3494]<=16'd4867; ROM2[3494]<=16'd0; ROM3[3494]<=16'd23842; ROM4[3494]<=16'd57335;
ROM1[3495]<=16'd4860; ROM2[3495]<=16'd0; ROM3[3495]<=16'd23853; ROM4[3495]<=16'd57344;
ROM1[3496]<=16'd4850; ROM2[3496]<=16'd0; ROM3[3496]<=16'd23859; ROM4[3496]<=16'd57348;
ROM1[3497]<=16'd4845; ROM2[3497]<=16'd0; ROM3[3497]<=16'd23849; ROM4[3497]<=16'd57341;
ROM1[3498]<=16'd4862; ROM2[3498]<=16'd0; ROM3[3498]<=16'd23838; ROM4[3498]<=16'd57335;
ROM1[3499]<=16'd4895; ROM2[3499]<=16'd0; ROM3[3499]<=16'd23831; ROM4[3499]<=16'd57339;
ROM1[3500]<=16'd4898; ROM2[3500]<=16'd0; ROM3[3500]<=16'd23831; ROM4[3500]<=16'd57337;
ROM1[3501]<=16'd4877; ROM2[3501]<=16'd0; ROM3[3501]<=16'd23830; ROM4[3501]<=16'd57330;
ROM1[3502]<=16'd4844; ROM2[3502]<=16'd0; ROM3[3502]<=16'd23824; ROM4[3502]<=16'd57317;
ROM1[3503]<=16'd4828; ROM2[3503]<=16'd0; ROM3[3503]<=16'd23829; ROM4[3503]<=16'd57313;
ROM1[3504]<=16'd4813; ROM2[3504]<=16'd0; ROM3[3504]<=16'd23832; ROM4[3504]<=16'd57313;
ROM1[3505]<=16'd4810; ROM2[3505]<=16'd0; ROM3[3505]<=16'd23831; ROM4[3505]<=16'd57310;
ROM1[3506]<=16'd4841; ROM2[3506]<=16'd0; ROM3[3506]<=16'd23835; ROM4[3506]<=16'd57321;
ROM1[3507]<=16'd4873; ROM2[3507]<=16'd0; ROM3[3507]<=16'd23825; ROM4[3507]<=16'd57321;
ROM1[3508]<=16'd4885; ROM2[3508]<=16'd0; ROM3[3508]<=16'd23822; ROM4[3508]<=16'd57320;
ROM1[3509]<=16'd4873; ROM2[3509]<=16'd0; ROM3[3509]<=16'd23828; ROM4[3509]<=16'd57326;
ROM1[3510]<=16'd4863; ROM2[3510]<=16'd0; ROM3[3510]<=16'd23848; ROM4[3510]<=16'd57336;
ROM1[3511]<=16'd4851; ROM2[3511]<=16'd0; ROM3[3511]<=16'd23850; ROM4[3511]<=16'd57332;
ROM1[3512]<=16'd4813; ROM2[3512]<=16'd0; ROM3[3512]<=16'd23825; ROM4[3512]<=16'd57305;
ROM1[3513]<=16'd4802; ROM2[3513]<=16'd0; ROM3[3513]<=16'd23819; ROM4[3513]<=16'd57297;
ROM1[3514]<=16'd4813; ROM2[3514]<=16'd0; ROM3[3514]<=16'd23810; ROM4[3514]<=16'd57293;
ROM1[3515]<=16'd4833; ROM2[3515]<=16'd0; ROM3[3515]<=16'd23792; ROM4[3515]<=16'd57285;
ROM1[3516]<=16'd4865; ROM2[3516]<=16'd0; ROM3[3516]<=16'd23794; ROM4[3516]<=16'd57296;
ROM1[3517]<=16'd4868; ROM2[3517]<=16'd0; ROM3[3517]<=16'd23802; ROM4[3517]<=16'd57307;
ROM1[3518]<=16'd4844; ROM2[3518]<=16'd0; ROM3[3518]<=16'd23801; ROM4[3518]<=16'd57301;
ROM1[3519]<=16'd4829; ROM2[3519]<=16'd0; ROM3[3519]<=16'd23812; ROM4[3519]<=16'd57300;
ROM1[3520]<=16'd4827; ROM2[3520]<=16'd0; ROM3[3520]<=16'd23831; ROM4[3520]<=16'd57313;
ROM1[3521]<=16'd4819; ROM2[3521]<=16'd0; ROM3[3521]<=16'd23841; ROM4[3521]<=16'd57322;
ROM1[3522]<=16'd4814; ROM2[3522]<=16'd0; ROM3[3522]<=16'd23832; ROM4[3522]<=16'd57314;
ROM1[3523]<=16'd4834; ROM2[3523]<=16'd0; ROM3[3523]<=16'd23819; ROM4[3523]<=16'd57309;
ROM1[3524]<=16'd4869; ROM2[3524]<=16'd0; ROM3[3524]<=16'd23808; ROM4[3524]<=16'd57310;
ROM1[3525]<=16'd4869; ROM2[3525]<=16'd0; ROM3[3525]<=16'd23801; ROM4[3525]<=16'd57303;
ROM1[3526]<=16'd4852; ROM2[3526]<=16'd0; ROM3[3526]<=16'd23801; ROM4[3526]<=16'd57300;
ROM1[3527]<=16'd4830; ROM2[3527]<=16'd0; ROM3[3527]<=16'd23806; ROM4[3527]<=16'd57300;
ROM1[3528]<=16'd4813; ROM2[3528]<=16'd0; ROM3[3528]<=16'd23809; ROM4[3528]<=16'd57298;
ROM1[3529]<=16'd4801; ROM2[3529]<=16'd0; ROM3[3529]<=16'd23816; ROM4[3529]<=16'd57298;
ROM1[3530]<=16'd4800; ROM2[3530]<=16'd0; ROM3[3530]<=16'd23818; ROM4[3530]<=16'd57298;
ROM1[3531]<=16'd4822; ROM2[3531]<=16'd0; ROM3[3531]<=16'd23814; ROM4[3531]<=16'd57303;
ROM1[3532]<=16'd4861; ROM2[3532]<=16'd0; ROM3[3532]<=16'd23809; ROM4[3532]<=16'd57311;
ROM1[3533]<=16'd4896; ROM2[3533]<=16'd0; ROM3[3533]<=16'd23819; ROM4[3533]<=16'd57326;
ROM1[3534]<=16'd4894; ROM2[3534]<=16'd0; ROM3[3534]<=16'd23834; ROM4[3534]<=16'd57340;
ROM1[3535]<=16'd4867; ROM2[3535]<=16'd0; ROM3[3535]<=16'd23833; ROM4[3535]<=16'd57334;
ROM1[3536]<=16'd4855; ROM2[3536]<=16'd0; ROM3[3536]<=16'd23842; ROM4[3536]<=16'd57333;
ROM1[3537]<=16'd4825; ROM2[3537]<=16'd0; ROM3[3537]<=16'd23832; ROM4[3537]<=16'd57320;
ROM1[3538]<=16'd4793; ROM2[3538]<=16'd0; ROM3[3538]<=16'd23807; ROM4[3538]<=16'd57295;
ROM1[3539]<=16'd4805; ROM2[3539]<=16'd0; ROM3[3539]<=16'd23806; ROM4[3539]<=16'd57298;
ROM1[3540]<=16'd4842; ROM2[3540]<=16'd0; ROM3[3540]<=16'd23806; ROM4[3540]<=16'd57306;
ROM1[3541]<=16'd4881; ROM2[3541]<=16'd0; ROM3[3541]<=16'd23813; ROM4[3541]<=16'd57324;
ROM1[3542]<=16'd4878; ROM2[3542]<=16'd0; ROM3[3542]<=16'd23819; ROM4[3542]<=16'd57327;
ROM1[3543]<=16'd4854; ROM2[3543]<=16'd0; ROM3[3543]<=16'd23820; ROM4[3543]<=16'd57317;
ROM1[3544]<=16'd4835; ROM2[3544]<=16'd0; ROM3[3544]<=16'd23825; ROM4[3544]<=16'd57315;
ROM1[3545]<=16'd4817; ROM2[3545]<=16'd0; ROM3[3545]<=16'd23828; ROM4[3545]<=16'd57312;
ROM1[3546]<=16'd4816; ROM2[3546]<=16'd0; ROM3[3546]<=16'd23842; ROM4[3546]<=16'd57324;
ROM1[3547]<=16'd4830; ROM2[3547]<=16'd0; ROM3[3547]<=16'd23847; ROM4[3547]<=16'd57330;
ROM1[3548]<=16'd4872; ROM2[3548]<=16'd0; ROM3[3548]<=16'd23851; ROM4[3548]<=16'd57343;
ROM1[3549]<=16'd4902; ROM2[3549]<=16'd0; ROM3[3549]<=16'd23833; ROM4[3549]<=16'd57337;
ROM1[3550]<=16'd4894; ROM2[3550]<=16'd0; ROM3[3550]<=16'd23815; ROM4[3550]<=16'd57323;
ROM1[3551]<=16'd4883; ROM2[3551]<=16'd0; ROM3[3551]<=16'd23826; ROM4[3551]<=16'd57329;
ROM1[3552]<=16'd4849; ROM2[3552]<=16'd0; ROM3[3552]<=16'd23815; ROM4[3552]<=16'd57315;
ROM1[3553]<=16'd4826; ROM2[3553]<=16'd0; ROM3[3553]<=16'd23807; ROM4[3553]<=16'd57303;
ROM1[3554]<=16'd4825; ROM2[3554]<=16'd0; ROM3[3554]<=16'd23825; ROM4[3554]<=16'd57317;
ROM1[3555]<=16'd4824; ROM2[3555]<=16'd0; ROM3[3555]<=16'd23821; ROM4[3555]<=16'd57317;
ROM1[3556]<=16'd4833; ROM2[3556]<=16'd0; ROM3[3556]<=16'd23804; ROM4[3556]<=16'd57307;
ROM1[3557]<=16'd4868; ROM2[3557]<=16'd0; ROM3[3557]<=16'd23794; ROM4[3557]<=16'd57311;
ROM1[3558]<=16'd4891; ROM2[3558]<=16'd0; ROM3[3558]<=16'd23798; ROM4[3558]<=16'd57320;
ROM1[3559]<=16'd4876; ROM2[3559]<=16'd0; ROM3[3559]<=16'd23803; ROM4[3559]<=16'd57319;
ROM1[3560]<=16'd4855; ROM2[3560]<=16'd0; ROM3[3560]<=16'd23806; ROM4[3560]<=16'd57316;
ROM1[3561]<=16'd4848; ROM2[3561]<=16'd0; ROM3[3561]<=16'd23817; ROM4[3561]<=16'd57323;
ROM1[3562]<=16'd4837; ROM2[3562]<=16'd0; ROM3[3562]<=16'd23829; ROM4[3562]<=16'd57327;
ROM1[3563]<=16'd4837; ROM2[3563]<=16'd0; ROM3[3563]<=16'd23840; ROM4[3563]<=16'd57334;
ROM1[3564]<=16'd4854; ROM2[3564]<=16'd0; ROM3[3564]<=16'd23847; ROM4[3564]<=16'd57344;
ROM1[3565]<=16'd4865; ROM2[3565]<=16'd0; ROM3[3565]<=16'd23829; ROM4[3565]<=16'd57329;
ROM1[3566]<=16'd4868; ROM2[3566]<=16'd0; ROM3[3566]<=16'd23805; ROM4[3566]<=16'd57307;
ROM1[3567]<=16'd4858; ROM2[3567]<=16'd0; ROM3[3567]<=16'd23803; ROM4[3567]<=16'd57303;
ROM1[3568]<=16'd4840; ROM2[3568]<=16'd0; ROM3[3568]<=16'd23813; ROM4[3568]<=16'd57302;
ROM1[3569]<=16'd4840; ROM2[3569]<=16'd0; ROM3[3569]<=16'd23838; ROM4[3569]<=16'd57318;
ROM1[3570]<=16'd4840; ROM2[3570]<=16'd0; ROM3[3570]<=16'd23850; ROM4[3570]<=16'd57328;
ROM1[3571]<=16'd4816; ROM2[3571]<=16'd0; ROM3[3571]<=16'd23840; ROM4[3571]<=16'd57316;
ROM1[3572]<=16'd4811; ROM2[3572]<=16'd0; ROM3[3572]<=16'd23830; ROM4[3572]<=16'd57306;
ROM1[3573]<=16'd4837; ROM2[3573]<=16'd0; ROM3[3573]<=16'd23821; ROM4[3573]<=16'd57307;
ROM1[3574]<=16'd4879; ROM2[3574]<=16'd0; ROM3[3574]<=16'd23821; ROM4[3574]<=16'd57324;
ROM1[3575]<=16'd4903; ROM2[3575]<=16'd0; ROM3[3575]<=16'd23838; ROM4[3575]<=16'd57344;
ROM1[3576]<=16'd4883; ROM2[3576]<=16'd0; ROM3[3576]<=16'd23840; ROM4[3576]<=16'd57338;
ROM1[3577]<=16'd4840; ROM2[3577]<=16'd0; ROM3[3577]<=16'd23834; ROM4[3577]<=16'd57323;
ROM1[3578]<=16'd4815; ROM2[3578]<=16'd0; ROM3[3578]<=16'd23834; ROM4[3578]<=16'd57313;
ROM1[3579]<=16'd4796; ROM2[3579]<=16'd0; ROM3[3579]<=16'd23833; ROM4[3579]<=16'd57310;
ROM1[3580]<=16'd4803; ROM2[3580]<=16'd0; ROM3[3580]<=16'd23838; ROM4[3580]<=16'd57316;
ROM1[3581]<=16'd4827; ROM2[3581]<=16'd0; ROM3[3581]<=16'd23830; ROM4[3581]<=16'd57318;
ROM1[3582]<=16'd4858; ROM2[3582]<=16'd0; ROM3[3582]<=16'd23816; ROM4[3582]<=16'd57317;
ROM1[3583]<=16'd4871; ROM2[3583]<=16'd0; ROM3[3583]<=16'd23811; ROM4[3583]<=16'd57319;
ROM1[3584]<=16'd4861; ROM2[3584]<=16'd0; ROM3[3584]<=16'd23819; ROM4[3584]<=16'd57322;
ROM1[3585]<=16'd4850; ROM2[3585]<=16'd0; ROM3[3585]<=16'd23830; ROM4[3585]<=16'd57328;
ROM1[3586]<=16'd4845; ROM2[3586]<=16'd0; ROM3[3586]<=16'd23840; ROM4[3586]<=16'd57332;
ROM1[3587]<=16'd4831; ROM2[3587]<=16'd0; ROM3[3587]<=16'd23839; ROM4[3587]<=16'd57325;
ROM1[3588]<=16'd4821; ROM2[3588]<=16'd0; ROM3[3588]<=16'd23837; ROM4[3588]<=16'd57322;
ROM1[3589]<=16'd4824; ROM2[3589]<=16'd0; ROM3[3589]<=16'd23828; ROM4[3589]<=16'd57313;
ROM1[3590]<=16'd4848; ROM2[3590]<=16'd0; ROM3[3590]<=16'd23810; ROM4[3590]<=16'd57305;
ROM1[3591]<=16'd4870; ROM2[3591]<=16'd0; ROM3[3591]<=16'd23794; ROM4[3591]<=16'd57301;
ROM1[3592]<=16'd4863; ROM2[3592]<=16'd0; ROM3[3592]<=16'd23792; ROM4[3592]<=16'd57294;
ROM1[3593]<=16'd4862; ROM2[3593]<=16'd0; ROM3[3593]<=16'd23811; ROM4[3593]<=16'd57306;
ROM1[3594]<=16'd4869; ROM2[3594]<=16'd0; ROM3[3594]<=16'd23841; ROM4[3594]<=16'd57325;
ROM1[3595]<=16'd4857; ROM2[3595]<=16'd0; ROM3[3595]<=16'd23846; ROM4[3595]<=16'd57322;
ROM1[3596]<=16'd4826; ROM2[3596]<=16'd0; ROM3[3596]<=16'd23826; ROM4[3596]<=16'd57298;
ROM1[3597]<=16'd4827; ROM2[3597]<=16'd0; ROM3[3597]<=16'd23816; ROM4[3597]<=16'd57292;
ROM1[3598]<=16'd4852; ROM2[3598]<=16'd0; ROM3[3598]<=16'd23809; ROM4[3598]<=16'd57293;
ROM1[3599]<=16'd4883; ROM2[3599]<=16'd0; ROM3[3599]<=16'd23799; ROM4[3599]<=16'd57293;
ROM1[3600]<=16'd4897; ROM2[3600]<=16'd0; ROM3[3600]<=16'd23807; ROM4[3600]<=16'd57307;
ROM1[3601]<=16'd4878; ROM2[3601]<=16'd0; ROM3[3601]<=16'd23817; ROM4[3601]<=16'd57310;
ROM1[3602]<=16'd4846; ROM2[3602]<=16'd0; ROM3[3602]<=16'd23817; ROM4[3602]<=16'd57304;
ROM1[3603]<=16'd4833; ROM2[3603]<=16'd0; ROM3[3603]<=16'd23830; ROM4[3603]<=16'd57308;
ROM1[3604]<=16'd4825; ROM2[3604]<=16'd0; ROM3[3604]<=16'd23849; ROM4[3604]<=16'd57317;
ROM1[3605]<=16'd4825; ROM2[3605]<=16'd0; ROM3[3605]<=16'd23852; ROM4[3605]<=16'd57316;
ROM1[3606]<=16'd4832; ROM2[3606]<=16'd0; ROM3[3606]<=16'd23832; ROM4[3606]<=16'd57300;
ROM1[3607]<=16'd4861; ROM2[3607]<=16'd0; ROM3[3607]<=16'd23815; ROM4[3607]<=16'd57297;
ROM1[3608]<=16'd4880; ROM2[3608]<=16'd0; ROM3[3608]<=16'd23818; ROM4[3608]<=16'd57306;
ROM1[3609]<=16'd4866; ROM2[3609]<=16'd0; ROM3[3609]<=16'd23826; ROM4[3609]<=16'd57313;
ROM1[3610]<=16'd4853; ROM2[3610]<=16'd0; ROM3[3610]<=16'd23837; ROM4[3610]<=16'd57315;
ROM1[3611]<=16'd4849; ROM2[3611]<=16'd0; ROM3[3611]<=16'd23852; ROM4[3611]<=16'd57321;
ROM1[3612]<=16'd4845; ROM2[3612]<=16'd0; ROM3[3612]<=16'd23861; ROM4[3612]<=16'd57329;
ROM1[3613]<=16'd4839; ROM2[3613]<=16'd0; ROM3[3613]<=16'd23860; ROM4[3613]<=16'd57329;
ROM1[3614]<=16'd4854; ROM2[3614]<=16'd0; ROM3[3614]<=16'd23860; ROM4[3614]<=16'd57334;
ROM1[3615]<=16'd4884; ROM2[3615]<=16'd0; ROM3[3615]<=16'd23849; ROM4[3615]<=16'd57339;
ROM1[3616]<=16'd4904; ROM2[3616]<=16'd0; ROM3[3616]<=16'd23838; ROM4[3616]<=16'd57338;
ROM1[3617]<=16'd4909; ROM2[3617]<=16'd0; ROM3[3617]<=16'd23851; ROM4[3617]<=16'd57351;
ROM1[3618]<=16'd4890; ROM2[3618]<=16'd0; ROM3[3618]<=16'd23859; ROM4[3618]<=16'd57353;
ROM1[3619]<=16'd4858; ROM2[3619]<=16'd0; ROM3[3619]<=16'd23855; ROM4[3619]<=16'd57342;
ROM1[3620]<=16'd4836; ROM2[3620]<=16'd0; ROM3[3620]<=16'd23853; ROM4[3620]<=16'd57337;
ROM1[3621]<=16'd4814; ROM2[3621]<=16'd0; ROM3[3621]<=16'd23844; ROM4[3621]<=16'd57322;
ROM1[3622]<=16'd4823; ROM2[3622]<=16'd0; ROM3[3622]<=16'd23843; ROM4[3622]<=16'd57323;
ROM1[3623]<=16'd4850; ROM2[3623]<=16'd0; ROM3[3623]<=16'd23841; ROM4[3623]<=16'd57325;
ROM1[3624]<=16'd4881; ROM2[3624]<=16'd0; ROM3[3624]<=16'd23831; ROM4[3624]<=16'd57323;
ROM1[3625]<=16'd4882; ROM2[3625]<=16'd0; ROM3[3625]<=16'd23824; ROM4[3625]<=16'd57319;
ROM1[3626]<=16'd4860; ROM2[3626]<=16'd0; ROM3[3626]<=16'd23823; ROM4[3626]<=16'd57313;
ROM1[3627]<=16'd4863; ROM2[3627]<=16'd0; ROM3[3627]<=16'd23848; ROM4[3627]<=16'd57332;
ROM1[3628]<=16'd4856; ROM2[3628]<=16'd0; ROM3[3628]<=16'd23856; ROM4[3628]<=16'd57338;
ROM1[3629]<=16'd4812; ROM2[3629]<=16'd0; ROM3[3629]<=16'd23835; ROM4[3629]<=16'd57305;
ROM1[3630]<=16'd4799; ROM2[3630]<=16'd0; ROM3[3630]<=16'd23826; ROM4[3630]<=16'd57292;
ROM1[3631]<=16'd4813; ROM2[3631]<=16'd0; ROM3[3631]<=16'd23811; ROM4[3631]<=16'd57285;
ROM1[3632]<=16'd4850; ROM2[3632]<=16'd0; ROM3[3632]<=16'd23799; ROM4[3632]<=16'd57283;
ROM1[3633]<=16'd4887; ROM2[3633]<=16'd0; ROM3[3633]<=16'd23804; ROM4[3633]<=16'd57301;
ROM1[3634]<=16'd4891; ROM2[3634]<=16'd0; ROM3[3634]<=16'd23818; ROM4[3634]<=16'd57314;
ROM1[3635]<=16'd4875; ROM2[3635]<=16'd0; ROM3[3635]<=16'd23830; ROM4[3635]<=16'd57318;
ROM1[3636]<=16'd4858; ROM2[3636]<=16'd0; ROM3[3636]<=16'd23833; ROM4[3636]<=16'd57316;
ROM1[3637]<=16'd4833; ROM2[3637]<=16'd0; ROM3[3637]<=16'd23834; ROM4[3637]<=16'd57311;
ROM1[3638]<=16'd4823; ROM2[3638]<=16'd0; ROM3[3638]<=16'd23832; ROM4[3638]<=16'd57309;
ROM1[3639]<=16'd4837; ROM2[3639]<=16'd0; ROM3[3639]<=16'd23824; ROM4[3639]<=16'd57306;
ROM1[3640]<=16'd4861; ROM2[3640]<=16'd0; ROM3[3640]<=16'd23806; ROM4[3640]<=16'd57300;
ROM1[3641]<=16'd4891; ROM2[3641]<=16'd0; ROM3[3641]<=16'd23804; ROM4[3641]<=16'd57307;
ROM1[3642]<=16'd4883; ROM2[3642]<=16'd0; ROM3[3642]<=16'd23806; ROM4[3642]<=16'd57306;
ROM1[3643]<=16'd4854; ROM2[3643]<=16'd0; ROM3[3643]<=16'd23802; ROM4[3643]<=16'd57294;
ROM1[3644]<=16'd4834; ROM2[3644]<=16'd0; ROM3[3644]<=16'd23809; ROM4[3644]<=16'd57291;
ROM1[3645]<=16'd4826; ROM2[3645]<=16'd0; ROM3[3645]<=16'd23817; ROM4[3645]<=16'd57294;
ROM1[3646]<=16'd4815; ROM2[3646]<=16'd0; ROM3[3646]<=16'd23819; ROM4[3646]<=16'd57292;
ROM1[3647]<=16'd4815; ROM2[3647]<=16'd0; ROM3[3647]<=16'd23808; ROM4[3647]<=16'd57285;
ROM1[3648]<=16'd4838; ROM2[3648]<=16'd0; ROM3[3648]<=16'd23797; ROM4[3648]<=16'd57279;
ROM1[3649]<=16'd4872; ROM2[3649]<=16'd0; ROM3[3649]<=16'd23790; ROM4[3649]<=16'd57280;
ROM1[3650]<=16'd4883; ROM2[3650]<=16'd0; ROM3[3650]<=16'd23791; ROM4[3650]<=16'd57285;
ROM1[3651]<=16'd4862; ROM2[3651]<=16'd0; ROM3[3651]<=16'd23793; ROM4[3651]<=16'd57281;
ROM1[3652]<=16'd4842; ROM2[3652]<=16'd0; ROM3[3652]<=16'd23795; ROM4[3652]<=16'd57278;
ROM1[3653]<=16'd4838; ROM2[3653]<=16'd0; ROM3[3653]<=16'd23808; ROM4[3653]<=16'd57287;
ROM1[3654]<=16'd4830; ROM2[3654]<=16'd0; ROM3[3654]<=16'd23816; ROM4[3654]<=16'd57290;
ROM1[3655]<=16'd4829; ROM2[3655]<=16'd0; ROM3[3655]<=16'd23816; ROM4[3655]<=16'd57288;
ROM1[3656]<=16'd4850; ROM2[3656]<=16'd0; ROM3[3656]<=16'd23813; ROM4[3656]<=16'd57292;
ROM1[3657]<=16'd4875; ROM2[3657]<=16'd0; ROM3[3657]<=16'd23794; ROM4[3657]<=16'd57289;
ROM1[3658]<=16'd4880; ROM2[3658]<=16'd0; ROM3[3658]<=16'd23787; ROM4[3658]<=16'd57284;
ROM1[3659]<=16'd4877; ROM2[3659]<=16'd0; ROM3[3659]<=16'd23797; ROM4[3659]<=16'd57293;
ROM1[3660]<=16'd4871; ROM2[3660]<=16'd0; ROM3[3660]<=16'd23812; ROM4[3660]<=16'd57308;
ROM1[3661]<=16'd4863; ROM2[3661]<=16'd0; ROM3[3661]<=16'd23819; ROM4[3661]<=16'd57305;
ROM1[3662]<=16'd4845; ROM2[3662]<=16'd0; ROM3[3662]<=16'd23816; ROM4[3662]<=16'd57297;
ROM1[3663]<=16'd4848; ROM2[3663]<=16'd0; ROM3[3663]<=16'd23829; ROM4[3663]<=16'd57311;
ROM1[3664]<=16'd4875; ROM2[3664]<=16'd0; ROM3[3664]<=16'd23840; ROM4[3664]<=16'd57329;
ROM1[3665]<=16'd4911; ROM2[3665]<=16'd0; ROM3[3665]<=16'd23834; ROM4[3665]<=16'd57336;
ROM1[3666]<=16'd4925; ROM2[3666]<=16'd0; ROM3[3666]<=16'd23813; ROM4[3666]<=16'd57325;
ROM1[3667]<=16'd4902; ROM2[3667]<=16'd0; ROM3[3667]<=16'd23800; ROM4[3667]<=16'd57310;
ROM1[3668]<=16'd4868; ROM2[3668]<=16'd0; ROM3[3668]<=16'd23796; ROM4[3668]<=16'd57299;
ROM1[3669]<=16'd4842; ROM2[3669]<=16'd0; ROM3[3669]<=16'd23797; ROM4[3669]<=16'd57295;
ROM1[3670]<=16'd4847; ROM2[3670]<=16'd0; ROM3[3670]<=16'd23822; ROM4[3670]<=16'd57315;
ROM1[3671]<=16'd4859; ROM2[3671]<=16'd0; ROM3[3671]<=16'd23848; ROM4[3671]<=16'd57334;
ROM1[3672]<=16'd4850; ROM2[3672]<=16'd0; ROM3[3672]<=16'd23834; ROM4[3672]<=16'd57321;
ROM1[3673]<=16'd4871; ROM2[3673]<=16'd0; ROM3[3673]<=16'd23823; ROM4[3673]<=16'd57317;
ROM1[3674]<=16'd4898; ROM2[3674]<=16'd0; ROM3[3674]<=16'd23809; ROM4[3674]<=16'd57317;
ROM1[3675]<=16'd4877; ROM2[3675]<=16'd0; ROM3[3675]<=16'd23787; ROM4[3675]<=16'd57301;
ROM1[3676]<=16'd4867; ROM2[3676]<=16'd0; ROM3[3676]<=16'd23805; ROM4[3676]<=16'd57305;
ROM1[3677]<=16'd4856; ROM2[3677]<=16'd0; ROM3[3677]<=16'd23826; ROM4[3677]<=16'd57316;
ROM1[3678]<=16'd4845; ROM2[3678]<=16'd0; ROM3[3678]<=16'd23838; ROM4[3678]<=16'd57320;
ROM1[3679]<=16'd4840; ROM2[3679]<=16'd0; ROM3[3679]<=16'd23852; ROM4[3679]<=16'd57327;
ROM1[3680]<=16'd4840; ROM2[3680]<=16'd0; ROM3[3680]<=16'd23852; ROM4[3680]<=16'd57329;
ROM1[3681]<=16'd4853; ROM2[3681]<=16'd0; ROM3[3681]<=16'd23841; ROM4[3681]<=16'd57322;
ROM1[3682]<=16'd4889; ROM2[3682]<=16'd0; ROM3[3682]<=16'd23837; ROM4[3682]<=16'd57328;
ROM1[3683]<=16'd4912; ROM2[3683]<=16'd0; ROM3[3683]<=16'd23838; ROM4[3683]<=16'd57334;
ROM1[3684]<=16'd4885; ROM2[3684]<=16'd0; ROM3[3684]<=16'd23829; ROM4[3684]<=16'd57317;
ROM1[3685]<=16'd4845; ROM2[3685]<=16'd0; ROM3[3685]<=16'd23821; ROM4[3685]<=16'd57302;
ROM1[3686]<=16'd4818; ROM2[3686]<=16'd0; ROM3[3686]<=16'd23817; ROM4[3686]<=16'd57292;
ROM1[3687]<=16'd4788; ROM2[3687]<=16'd0; ROM3[3687]<=16'd23809; ROM4[3687]<=16'd57274;
ROM1[3688]<=16'd4782; ROM2[3688]<=16'd0; ROM3[3688]<=16'd23804; ROM4[3688]<=16'd57271;
ROM1[3689]<=16'd4802; ROM2[3689]<=16'd0; ROM3[3689]<=16'd23799; ROM4[3689]<=16'd57277;
ROM1[3690]<=16'd4830; ROM2[3690]<=16'd0; ROM3[3690]<=16'd23786; ROM4[3690]<=16'd57275;
ROM1[3691]<=16'd4857; ROM2[3691]<=16'd0; ROM3[3691]<=16'd23782; ROM4[3691]<=16'd57282;
ROM1[3692]<=16'd4856; ROM2[3692]<=16'd0; ROM3[3692]<=16'd23789; ROM4[3692]<=16'd57292;
ROM1[3693]<=16'd4839; ROM2[3693]<=16'd0; ROM3[3693]<=16'd23793; ROM4[3693]<=16'd57291;
ROM1[3694]<=16'd4822; ROM2[3694]<=16'd0; ROM3[3694]<=16'd23797; ROM4[3694]<=16'd57287;
ROM1[3695]<=16'd4808; ROM2[3695]<=16'd0; ROM3[3695]<=16'd23795; ROM4[3695]<=16'd57285;
ROM1[3696]<=16'd4805; ROM2[3696]<=16'd0; ROM3[3696]<=16'd23800; ROM4[3696]<=16'd57290;
ROM1[3697]<=16'd4819; ROM2[3697]<=16'd0; ROM3[3697]<=16'd23802; ROM4[3697]<=16'd57294;
ROM1[3698]<=16'd4850; ROM2[3698]<=16'd0; ROM3[3698]<=16'd23793; ROM4[3698]<=16'd57299;
ROM1[3699]<=16'd4881; ROM2[3699]<=16'd0; ROM3[3699]<=16'd23779; ROM4[3699]<=16'd57298;
ROM1[3700]<=16'd4887; ROM2[3700]<=16'd0; ROM3[3700]<=16'd23783; ROM4[3700]<=16'd57299;
ROM1[3701]<=16'd4891; ROM2[3701]<=16'd0; ROM3[3701]<=16'd23809; ROM4[3701]<=16'd57318;
ROM1[3702]<=16'd4873; ROM2[3702]<=16'd0; ROM3[3702]<=16'd23810; ROM4[3702]<=16'd57315;
ROM1[3703]<=16'd4846; ROM2[3703]<=16'd0; ROM3[3703]<=16'd23800; ROM4[3703]<=16'd57299;
ROM1[3704]<=16'd4825; ROM2[3704]<=16'd0; ROM3[3704]<=16'd23800; ROM4[3704]<=16'd57296;
ROM1[3705]<=16'd4818; ROM2[3705]<=16'd0; ROM3[3705]<=16'd23791; ROM4[3705]<=16'd57292;
ROM1[3706]<=16'd4838; ROM2[3706]<=16'd0; ROM3[3706]<=16'd23783; ROM4[3706]<=16'd57288;
ROM1[3707]<=16'd4883; ROM2[3707]<=16'd0; ROM3[3707]<=16'd23781; ROM4[3707]<=16'd57297;
ROM1[3708]<=16'd4906; ROM2[3708]<=16'd0; ROM3[3708]<=16'd23784; ROM4[3708]<=16'd57308;
ROM1[3709]<=16'd4895; ROM2[3709]<=16'd0; ROM3[3709]<=16'd23795; ROM4[3709]<=16'd57310;
ROM1[3710]<=16'd4866; ROM2[3710]<=16'd0; ROM3[3710]<=16'd23797; ROM4[3710]<=16'd57303;
ROM1[3711]<=16'd4849; ROM2[3711]<=16'd0; ROM3[3711]<=16'd23807; ROM4[3711]<=16'd57306;
ROM1[3712]<=16'd4841; ROM2[3712]<=16'd0; ROM3[3712]<=16'd23820; ROM4[3712]<=16'd57309;
ROM1[3713]<=16'd4833; ROM2[3713]<=16'd0; ROM3[3713]<=16'd23813; ROM4[3713]<=16'd57298;
ROM1[3714]<=16'd4858; ROM2[3714]<=16'd0; ROM3[3714]<=16'd23819; ROM4[3714]<=16'd57305;
ROM1[3715]<=16'd4900; ROM2[3715]<=16'd0; ROM3[3715]<=16'd23821; ROM4[3715]<=16'd57320;
ROM1[3716]<=16'd4904; ROM2[3716]<=16'd0; ROM3[3716]<=16'd23792; ROM4[3716]<=16'd57300;
ROM1[3717]<=16'd4890; ROM2[3717]<=16'd0; ROM3[3717]<=16'd23788; ROM4[3717]<=16'd57295;
ROM1[3718]<=16'd4886; ROM2[3718]<=16'd0; ROM3[3718]<=16'd23810; ROM4[3718]<=16'd57317;
ROM1[3719]<=16'd4864; ROM2[3719]<=16'd0; ROM3[3719]<=16'd23813; ROM4[3719]<=16'd57312;
ROM1[3720]<=16'd4852; ROM2[3720]<=16'd0; ROM3[3720]<=16'd23820; ROM4[3720]<=16'd57312;
ROM1[3721]<=16'd4837; ROM2[3721]<=16'd0; ROM3[3721]<=16'd23828; ROM4[3721]<=16'd57312;
ROM1[3722]<=16'd4829; ROM2[3722]<=16'd0; ROM3[3722]<=16'd23814; ROM4[3722]<=16'd57301;
ROM1[3723]<=16'd4858; ROM2[3723]<=16'd0; ROM3[3723]<=16'd23808; ROM4[3723]<=16'd57303;
ROM1[3724]<=16'd4891; ROM2[3724]<=16'd0; ROM3[3724]<=16'd23805; ROM4[3724]<=16'd57306;
ROM1[3725]<=16'd4891; ROM2[3725]<=16'd0; ROM3[3725]<=16'd23801; ROM4[3725]<=16'd57304;
ROM1[3726]<=16'd4884; ROM2[3726]<=16'd0; ROM3[3726]<=16'd23819; ROM4[3726]<=16'd57313;
ROM1[3727]<=16'd4880; ROM2[3727]<=16'd0; ROM3[3727]<=16'd23842; ROM4[3727]<=16'd57325;
ROM1[3728]<=16'd4868; ROM2[3728]<=16'd0; ROM3[3728]<=16'd23844; ROM4[3728]<=16'd57329;
ROM1[3729]<=16'd4835; ROM2[3729]<=16'd0; ROM3[3729]<=16'd23834; ROM4[3729]<=16'd57311;
ROM1[3730]<=16'd4822; ROM2[3730]<=16'd0; ROM3[3730]<=16'd23823; ROM4[3730]<=16'd57298;
ROM1[3731]<=16'd4828; ROM2[3731]<=16'd0; ROM3[3731]<=16'd23803; ROM4[3731]<=16'd57289;
ROM1[3732]<=16'd4863; ROM2[3732]<=16'd0; ROM3[3732]<=16'd23793; ROM4[3732]<=16'd57286;
ROM1[3733]<=16'd4887; ROM2[3733]<=16'd0; ROM3[3733]<=16'd23794; ROM4[3733]<=16'd57298;
ROM1[3734]<=16'd4873; ROM2[3734]<=16'd0; ROM3[3734]<=16'd23795; ROM4[3734]<=16'd57296;
ROM1[3735]<=16'd4852; ROM2[3735]<=16'd0; ROM3[3735]<=16'd23801; ROM4[3735]<=16'd57292;
ROM1[3736]<=16'd4856; ROM2[3736]<=16'd0; ROM3[3736]<=16'd23825; ROM4[3736]<=16'd57310;
ROM1[3737]<=16'd4855; ROM2[3737]<=16'd0; ROM3[3737]<=16'd23844; ROM4[3737]<=16'd57323;
ROM1[3738]<=16'd4842; ROM2[3738]<=16'd0; ROM3[3738]<=16'd23834; ROM4[3738]<=16'd57313;
ROM1[3739]<=16'd4853; ROM2[3739]<=16'd0; ROM3[3739]<=16'd23824; ROM4[3739]<=16'd57307;
ROM1[3740]<=16'd4876; ROM2[3740]<=16'd0; ROM3[3740]<=16'd23805; ROM4[3740]<=16'd57298;
ROM1[3741]<=16'd4896; ROM2[3741]<=16'd0; ROM3[3741]<=16'd23791; ROM4[3741]<=16'd57298;
ROM1[3742]<=16'd4894; ROM2[3742]<=16'd0; ROM3[3742]<=16'd23798; ROM4[3742]<=16'd57303;
ROM1[3743]<=16'd4873; ROM2[3743]<=16'd0; ROM3[3743]<=16'd23800; ROM4[3743]<=16'd57298;
ROM1[3744]<=16'd4851; ROM2[3744]<=16'd0; ROM3[3744]<=16'd23801; ROM4[3744]<=16'd57296;
ROM1[3745]<=16'd4851; ROM2[3745]<=16'd0; ROM3[3745]<=16'd23818; ROM4[3745]<=16'd57307;
ROM1[3746]<=16'd4848; ROM2[3746]<=16'd0; ROM3[3746]<=16'd23832; ROM4[3746]<=16'd57319;
ROM1[3747]<=16'd4837; ROM2[3747]<=16'd0; ROM3[3747]<=16'd23818; ROM4[3747]<=16'd57306;
ROM1[3748]<=16'd4849; ROM2[3748]<=16'd0; ROM3[3748]<=16'd23796; ROM4[3748]<=16'd57292;
ROM1[3749]<=16'd4882; ROM2[3749]<=16'd0; ROM3[3749]<=16'd23788; ROM4[3749]<=16'd57297;
ROM1[3750]<=16'd4886; ROM2[3750]<=16'd0; ROM3[3750]<=16'd23789; ROM4[3750]<=16'd57303;
ROM1[3751]<=16'd4860; ROM2[3751]<=16'd0; ROM3[3751]<=16'd23783; ROM4[3751]<=16'd57293;
ROM1[3752]<=16'd4824; ROM2[3752]<=16'd0; ROM3[3752]<=16'd23780; ROM4[3752]<=16'd57284;
ROM1[3753]<=16'd4802; ROM2[3753]<=16'd0; ROM3[3753]<=16'd23780; ROM4[3753]<=16'd57278;
ROM1[3754]<=16'd4783; ROM2[3754]<=16'd0; ROM3[3754]<=16'd23780; ROM4[3754]<=16'd57271;
ROM1[3755]<=16'd4798; ROM2[3755]<=16'd0; ROM3[3755]<=16'd23797; ROM4[3755]<=16'd57287;
ROM1[3756]<=16'd4828; ROM2[3756]<=16'd0; ROM3[3756]<=16'd23802; ROM4[3756]<=16'd57300;
ROM1[3757]<=16'd4855; ROM2[3757]<=16'd0; ROM3[3757]<=16'd23785; ROM4[3757]<=16'd57296;
ROM1[3758]<=16'd4867; ROM2[3758]<=16'd0; ROM3[3758]<=16'd23778; ROM4[3758]<=16'd57293;
ROM1[3759]<=16'd4865; ROM2[3759]<=16'd0; ROM3[3759]<=16'd23792; ROM4[3759]<=16'd57305;
ROM1[3760]<=16'd4854; ROM2[3760]<=16'd0; ROM3[3760]<=16'd23806; ROM4[3760]<=16'd57309;
ROM1[3761]<=16'd4840; ROM2[3761]<=16'd0; ROM3[3761]<=16'd23809; ROM4[3761]<=16'd57305;
ROM1[3762]<=16'd4824; ROM2[3762]<=16'd0; ROM3[3762]<=16'd23813; ROM4[3762]<=16'd57304;
ROM1[3763]<=16'd4822; ROM2[3763]<=16'd0; ROM3[3763]<=16'd23824; ROM4[3763]<=16'd57308;
ROM1[3764]<=16'd4833; ROM2[3764]<=16'd0; ROM3[3764]<=16'd23819; ROM4[3764]<=16'd57305;
ROM1[3765]<=16'd4858; ROM2[3765]<=16'd0; ROM3[3765]<=16'd23800; ROM4[3765]<=16'd57301;
ROM1[3766]<=16'd4878; ROM2[3766]<=16'd0; ROM3[3766]<=16'd23784; ROM4[3766]<=16'd57296;
ROM1[3767]<=16'd4876; ROM2[3767]<=16'd0; ROM3[3767]<=16'd23785; ROM4[3767]<=16'd57293;
ROM1[3768]<=16'd4872; ROM2[3768]<=16'd0; ROM3[3768]<=16'd23803; ROM4[3768]<=16'd57307;
ROM1[3769]<=16'd4863; ROM2[3769]<=16'd0; ROM3[3769]<=16'd23822; ROM4[3769]<=16'd57316;
ROM1[3770]<=16'd4869; ROM2[3770]<=16'd0; ROM3[3770]<=16'd23847; ROM4[3770]<=16'd57334;
ROM1[3771]<=16'd4869; ROM2[3771]<=16'd0; ROM3[3771]<=16'd23858; ROM4[3771]<=16'd57344;
ROM1[3772]<=16'd4861; ROM2[3772]<=16'd0; ROM3[3772]<=16'd23841; ROM4[3772]<=16'd57325;
ROM1[3773]<=16'd4865; ROM2[3773]<=16'd0; ROM3[3773]<=16'd23814; ROM4[3773]<=16'd57304;
ROM1[3774]<=16'd4881; ROM2[3774]<=16'd0; ROM3[3774]<=16'd23792; ROM4[3774]<=16'd57290;
ROM1[3775]<=16'd4879; ROM2[3775]<=16'd0; ROM3[3775]<=16'd23787; ROM4[3775]<=16'd57288;
ROM1[3776]<=16'd4863; ROM2[3776]<=16'd0; ROM3[3776]<=16'd23793; ROM4[3776]<=16'd57290;
ROM1[3777]<=16'd4861; ROM2[3777]<=16'd0; ROM3[3777]<=16'd23814; ROM4[3777]<=16'd57304;
ROM1[3778]<=16'd4852; ROM2[3778]<=16'd0; ROM3[3778]<=16'd23825; ROM4[3778]<=16'd57310;
ROM1[3779]<=16'd4826; ROM2[3779]<=16'd0; ROM3[3779]<=16'd23818; ROM4[3779]<=16'd57299;
ROM1[3780]<=16'd4833; ROM2[3780]<=16'd0; ROM3[3780]<=16'd23820; ROM4[3780]<=16'd57304;
ROM1[3781]<=16'd4864; ROM2[3781]<=16'd0; ROM3[3781]<=16'd23816; ROM4[3781]<=16'd57310;
ROM1[3782]<=16'd4890; ROM2[3782]<=16'd0; ROM3[3782]<=16'd23795; ROM4[3782]<=16'd57303;
ROM1[3783]<=16'd4899; ROM2[3783]<=16'd0; ROM3[3783]<=16'd23789; ROM4[3783]<=16'd57305;
ROM1[3784]<=16'd4885; ROM2[3784]<=16'd0; ROM3[3784]<=16'd23797; ROM4[3784]<=16'd57310;
ROM1[3785]<=16'd4863; ROM2[3785]<=16'd0; ROM3[3785]<=16'd23800; ROM4[3785]<=16'd57307;
ROM1[3786]<=16'd4851; ROM2[3786]<=16'd0; ROM3[3786]<=16'd23800; ROM4[3786]<=16'd57303;
ROM1[3787]<=16'd4844; ROM2[3787]<=16'd0; ROM3[3787]<=16'd23804; ROM4[3787]<=16'd57302;
ROM1[3788]<=16'd4850; ROM2[3788]<=16'd0; ROM3[3788]<=16'd23811; ROM4[3788]<=16'd57304;
ROM1[3789]<=16'd4866; ROM2[3789]<=16'd0; ROM3[3789]<=16'd23820; ROM4[3789]<=16'd57311;
ROM1[3790]<=16'd4889; ROM2[3790]<=16'd0; ROM3[3790]<=16'd23811; ROM4[3790]<=16'd57309;
ROM1[3791]<=16'd4915; ROM2[3791]<=16'd0; ROM3[3791]<=16'd23805; ROM4[3791]<=16'd57313;
ROM1[3792]<=16'd4919; ROM2[3792]<=16'd0; ROM3[3792]<=16'd23818; ROM4[3792]<=16'd57327;
ROM1[3793]<=16'd4889; ROM2[3793]<=16'd0; ROM3[3793]<=16'd23813; ROM4[3793]<=16'd57312;
ROM1[3794]<=16'd4847; ROM2[3794]<=16'd0; ROM3[3794]<=16'd23796; ROM4[3794]<=16'd57287;
ROM1[3795]<=16'd4828; ROM2[3795]<=16'd0; ROM3[3795]<=16'd23801; ROM4[3795]<=16'd57283;
ROM1[3796]<=16'd4811; ROM2[3796]<=16'd0; ROM3[3796]<=16'd23797; ROM4[3796]<=16'd57273;
ROM1[3797]<=16'd4812; ROM2[3797]<=16'd0; ROM3[3797]<=16'd23785; ROM4[3797]<=16'd57265;
ROM1[3798]<=16'd4847; ROM2[3798]<=16'd0; ROM3[3798]<=16'd23785; ROM4[3798]<=16'd57275;
ROM1[3799]<=16'd4875; ROM2[3799]<=16'd0; ROM3[3799]<=16'd23770; ROM4[3799]<=16'd57276;
ROM1[3800]<=16'd4871; ROM2[3800]<=16'd0; ROM3[3800]<=16'd23766; ROM4[3800]<=16'd57271;
ROM1[3801]<=16'd4860; ROM2[3801]<=16'd0; ROM3[3801]<=16'd23780; ROM4[3801]<=16'd57279;
ROM1[3802]<=16'd4849; ROM2[3802]<=16'd0; ROM3[3802]<=16'd23795; ROM4[3802]<=16'd57289;
ROM1[3803]<=16'd4830; ROM2[3803]<=16'd0; ROM3[3803]<=16'd23792; ROM4[3803]<=16'd57284;
ROM1[3804]<=16'd4806; ROM2[3804]<=16'd0; ROM3[3804]<=16'd23785; ROM4[3804]<=16'd57274;
ROM1[3805]<=16'd4805; ROM2[3805]<=16'd0; ROM3[3805]<=16'd23783; ROM4[3805]<=16'd57273;
ROM1[3806]<=16'd4819; ROM2[3806]<=16'd0; ROM3[3806]<=16'd23770; ROM4[3806]<=16'd57269;
ROM1[3807]<=16'd4849; ROM2[3807]<=16'd0; ROM3[3807]<=16'd23760; ROM4[3807]<=16'd57268;
ROM1[3808]<=16'd4867; ROM2[3808]<=16'd0; ROM3[3808]<=16'd23764; ROM4[3808]<=16'd57276;
ROM1[3809]<=16'd4863; ROM2[3809]<=16'd0; ROM3[3809]<=16'd23774; ROM4[3809]<=16'd57281;
ROM1[3810]<=16'd4861; ROM2[3810]<=16'd0; ROM3[3810]<=16'd23800; ROM4[3810]<=16'd57299;
ROM1[3811]<=16'd4848; ROM2[3811]<=16'd0; ROM3[3811]<=16'd23805; ROM4[3811]<=16'd57301;
ROM1[3812]<=16'd4808; ROM2[3812]<=16'd0; ROM3[3812]<=16'd23784; ROM4[3812]<=16'd57279;
ROM1[3813]<=16'd4800; ROM2[3813]<=16'd0; ROM3[3813]<=16'd23786; ROM4[3813]<=16'd57280;
ROM1[3814]<=16'd4821; ROM2[3814]<=16'd0; ROM3[3814]<=16'd23789; ROM4[3814]<=16'd57288;
ROM1[3815]<=16'd4856; ROM2[3815]<=16'd0; ROM3[3815]<=16'd23779; ROM4[3815]<=16'd57290;
ROM1[3816]<=16'd4892; ROM2[3816]<=16'd0; ROM3[3816]<=16'd23784; ROM4[3816]<=16'd57303;
ROM1[3817]<=16'd4883; ROM2[3817]<=16'd0; ROM3[3817]<=16'd23785; ROM4[3817]<=16'd57302;
ROM1[3818]<=16'd4862; ROM2[3818]<=16'd0; ROM3[3818]<=16'd23784; ROM4[3818]<=16'd57297;
ROM1[3819]<=16'd4854; ROM2[3819]<=16'd0; ROM3[3819]<=16'd23798; ROM4[3819]<=16'd57303;
ROM1[3820]<=16'd4845; ROM2[3820]<=16'd0; ROM3[3820]<=16'd23806; ROM4[3820]<=16'd57306;
ROM1[3821]<=16'd4832; ROM2[3821]<=16'd0; ROM3[3821]<=16'd23807; ROM4[3821]<=16'd57299;
ROM1[3822]<=16'd4831; ROM2[3822]<=16'd0; ROM3[3822]<=16'd23797; ROM4[3822]<=16'd57289;
ROM1[3823]<=16'd4854; ROM2[3823]<=16'd0; ROM3[3823]<=16'd23788; ROM4[3823]<=16'd57292;
ROM1[3824]<=16'd4888; ROM2[3824]<=16'd0; ROM3[3824]<=16'd23784; ROM4[3824]<=16'd57296;
ROM1[3825]<=16'd4875; ROM2[3825]<=16'd0; ROM3[3825]<=16'd23769; ROM4[3825]<=16'd57284;
ROM1[3826]<=16'd4857; ROM2[3826]<=16'd0; ROM3[3826]<=16'd23773; ROM4[3826]<=16'd57283;
ROM1[3827]<=16'd4838; ROM2[3827]<=16'd0; ROM3[3827]<=16'd23780; ROM4[3827]<=16'd57282;
ROM1[3828]<=16'd4820; ROM2[3828]<=16'd0; ROM3[3828]<=16'd23786; ROM4[3828]<=16'd57282;
ROM1[3829]<=16'd4814; ROM2[3829]<=16'd0; ROM3[3829]<=16'd23798; ROM4[3829]<=16'd57288;
ROM1[3830]<=16'd4816; ROM2[3830]<=16'd0; ROM3[3830]<=16'd23799; ROM4[3830]<=16'd57289;
ROM1[3831]<=16'd4840; ROM2[3831]<=16'd0; ROM3[3831]<=16'd23795; ROM4[3831]<=16'd57287;
ROM1[3832]<=16'd4871; ROM2[3832]<=16'd0; ROM3[3832]<=16'd23777; ROM4[3832]<=16'd57280;
ROM1[3833]<=16'd4889; ROM2[3833]<=16'd0; ROM3[3833]<=16'd23775; ROM4[3833]<=16'd57288;
ROM1[3834]<=16'd4871; ROM2[3834]<=16'd0; ROM3[3834]<=16'd23785; ROM4[3834]<=16'd57290;
ROM1[3835]<=16'd4842; ROM2[3835]<=16'd0; ROM3[3835]<=16'd23786; ROM4[3835]<=16'd57283;
ROM1[3836]<=16'd4844; ROM2[3836]<=16'd0; ROM3[3836]<=16'd23803; ROM4[3836]<=16'd57295;
ROM1[3837]<=16'd4831; ROM2[3837]<=16'd0; ROM3[3837]<=16'd23812; ROM4[3837]<=16'd57299;
ROM1[3838]<=16'd4811; ROM2[3838]<=16'd0; ROM3[3838]<=16'd23797; ROM4[3838]<=16'd57285;
ROM1[3839]<=16'd4836; ROM2[3839]<=16'd0; ROM3[3839]<=16'd23809; ROM4[3839]<=16'd57296;
ROM1[3840]<=16'd4862; ROM2[3840]<=16'd0; ROM3[3840]<=16'd23801; ROM4[3840]<=16'd57296;
ROM1[3841]<=16'd4861; ROM2[3841]<=16'd0; ROM3[3841]<=16'd23768; ROM4[3841]<=16'd57273;
ROM1[3842]<=16'd4863; ROM2[3842]<=16'd0; ROM3[3842]<=16'd23778; ROM4[3842]<=16'd57282;
ROM1[3843]<=16'd4845; ROM2[3843]<=16'd0; ROM3[3843]<=16'd23784; ROM4[3843]<=16'd57284;
ROM1[3844]<=16'd4821; ROM2[3844]<=16'd0; ROM3[3844]<=16'd23783; ROM4[3844]<=16'd57277;
ROM1[3845]<=16'd4818; ROM2[3845]<=16'd0; ROM3[3845]<=16'd23797; ROM4[3845]<=16'd57289;
ROM1[3846]<=16'd4810; ROM2[3846]<=16'd0; ROM3[3846]<=16'd23804; ROM4[3846]<=16'd57292;
ROM1[3847]<=16'd4815; ROM2[3847]<=16'd0; ROM3[3847]<=16'd23800; ROM4[3847]<=16'd57289;
ROM1[3848]<=16'd4845; ROM2[3848]<=16'd0; ROM3[3848]<=16'd23790; ROM4[3848]<=16'd57291;
ROM1[3849]<=16'd4886; ROM2[3849]<=16'd0; ROM3[3849]<=16'd23791; ROM4[3849]<=16'd57302;
ROM1[3850]<=16'd4894; ROM2[3850]<=16'd0; ROM3[3850]<=16'd23791; ROM4[3850]<=16'd57304;
ROM1[3851]<=16'd4878; ROM2[3851]<=16'd0; ROM3[3851]<=16'd23793; ROM4[3851]<=16'd57302;
ROM1[3852]<=16'd4856; ROM2[3852]<=16'd0; ROM3[3852]<=16'd23801; ROM4[3852]<=16'd57296;
ROM1[3853]<=16'd4842; ROM2[3853]<=16'd0; ROM3[3853]<=16'd23804; ROM4[3853]<=16'd57290;
ROM1[3854]<=16'd4822; ROM2[3854]<=16'd0; ROM3[3854]<=16'd23804; ROM4[3854]<=16'd57286;
ROM1[3855]<=16'd4815; ROM2[3855]<=16'd0; ROM3[3855]<=16'd23799; ROM4[3855]<=16'd57283;
ROM1[3856]<=16'd4843; ROM2[3856]<=16'd0; ROM3[3856]<=16'd23796; ROM4[3856]<=16'd57289;
ROM1[3857]<=16'd4880; ROM2[3857]<=16'd0; ROM3[3857]<=16'd23790; ROM4[3857]<=16'd57296;
ROM1[3858]<=16'd4892; ROM2[3858]<=16'd0; ROM3[3858]<=16'd23784; ROM4[3858]<=16'd57293;
ROM1[3859]<=16'd4881; ROM2[3859]<=16'd0; ROM3[3859]<=16'd23790; ROM4[3859]<=16'd57293;
ROM1[3860]<=16'd4866; ROM2[3860]<=16'd0; ROM3[3860]<=16'd23803; ROM4[3860]<=16'd57302;
ROM1[3861]<=16'd4855; ROM2[3861]<=16'd0; ROM3[3861]<=16'd23808; ROM4[3861]<=16'd57304;
ROM1[3862]<=16'd4843; ROM2[3862]<=16'd0; ROM3[3862]<=16'd23816; ROM4[3862]<=16'd57307;
ROM1[3863]<=16'd4835; ROM2[3863]<=16'd0; ROM3[3863]<=16'd23817; ROM4[3863]<=16'd57307;
ROM1[3864]<=16'd4839; ROM2[3864]<=16'd0; ROM3[3864]<=16'd23807; ROM4[3864]<=16'd57301;
ROM1[3865]<=16'd4868; ROM2[3865]<=16'd0; ROM3[3865]<=16'd23800; ROM4[3865]<=16'd57305;
ROM1[3866]<=16'd4915; ROM2[3866]<=16'd0; ROM3[3866]<=16'd23813; ROM4[3866]<=16'd57326;
ROM1[3867]<=16'd4913; ROM2[3867]<=16'd0; ROM3[3867]<=16'd23815; ROM4[3867]<=16'd57328;
ROM1[3868]<=16'd4872; ROM2[3868]<=16'd0; ROM3[3868]<=16'd23796; ROM4[3868]<=16'd57300;
ROM1[3869]<=16'd4850; ROM2[3869]<=16'd0; ROM3[3869]<=16'd23796; ROM4[3869]<=16'd57292;
ROM1[3870]<=16'd4830; ROM2[3870]<=16'd0; ROM3[3870]<=16'd23797; ROM4[3870]<=16'd57286;
ROM1[3871]<=16'd4814; ROM2[3871]<=16'd0; ROM3[3871]<=16'd23795; ROM4[3871]<=16'd57280;
ROM1[3872]<=16'd4837; ROM2[3872]<=16'd0; ROM3[3872]<=16'd23805; ROM4[3872]<=16'd57293;
ROM1[3873]<=16'd4878; ROM2[3873]<=16'd0; ROM3[3873]<=16'd23812; ROM4[3873]<=16'd57307;
ROM1[3874]<=16'd4909; ROM2[3874]<=16'd0; ROM3[3874]<=16'd23800; ROM4[3874]<=16'd57304;
ROM1[3875]<=16'd4913; ROM2[3875]<=16'd0; ROM3[3875]<=16'd23799; ROM4[3875]<=16'd57304;
ROM1[3876]<=16'd4893; ROM2[3876]<=16'd0; ROM3[3876]<=16'd23812; ROM4[3876]<=16'd57308;
ROM1[3877]<=16'd4866; ROM2[3877]<=16'd0; ROM3[3877]<=16'd23813; ROM4[3877]<=16'd57300;
ROM1[3878]<=16'd4849; ROM2[3878]<=16'd0; ROM3[3878]<=16'd23817; ROM4[3878]<=16'd57299;
ROM1[3879]<=16'd4845; ROM2[3879]<=16'd0; ROM3[3879]<=16'd23828; ROM4[3879]<=16'd57308;
ROM1[3880]<=16'd4863; ROM2[3880]<=16'd0; ROM3[3880]<=16'd23834; ROM4[3880]<=16'd57323;
ROM1[3881]<=16'd4881; ROM2[3881]<=16'd0; ROM3[3881]<=16'd23820; ROM4[3881]<=16'd57322;
ROM1[3882]<=16'd4900; ROM2[3882]<=16'd0; ROM3[3882]<=16'd23796; ROM4[3882]<=16'd57310;
ROM1[3883]<=16'd4912; ROM2[3883]<=16'd0; ROM3[3883]<=16'd23791; ROM4[3883]<=16'd57310;
ROM1[3884]<=16'd4907; ROM2[3884]<=16'd0; ROM3[3884]<=16'd23803; ROM4[3884]<=16'd57318;
ROM1[3885]<=16'd4881; ROM2[3885]<=16'd0; ROM3[3885]<=16'd23806; ROM4[3885]<=16'd57311;
ROM1[3886]<=16'd4864; ROM2[3886]<=16'd0; ROM3[3886]<=16'd23813; ROM4[3886]<=16'd57314;
ROM1[3887]<=16'd4856; ROM2[3887]<=16'd0; ROM3[3887]<=16'd23829; ROM4[3887]<=16'd57328;
ROM1[3888]<=16'd4864; ROM2[3888]<=16'd0; ROM3[3888]<=16'd23845; ROM4[3888]<=16'd57341;
ROM1[3889]<=16'd4877; ROM2[3889]<=16'd0; ROM3[3889]<=16'd23839; ROM4[3889]<=16'd57340;
ROM1[3890]<=16'd4891; ROM2[3890]<=16'd0; ROM3[3890]<=16'd23813; ROM4[3890]<=16'd57319;
ROM1[3891]<=16'd4897; ROM2[3891]<=16'd0; ROM3[3891]<=16'd23787; ROM4[3891]<=16'd57302;
ROM1[3892]<=16'd4881; ROM2[3892]<=16'd0; ROM3[3892]<=16'd23786; ROM4[3892]<=16'd57297;
ROM1[3893]<=16'd4879; ROM2[3893]<=16'd0; ROM3[3893]<=16'd23809; ROM4[3893]<=16'd57315;
ROM1[3894]<=16'd4875; ROM2[3894]<=16'd0; ROM3[3894]<=16'd23830; ROM4[3894]<=16'd57328;
ROM1[3895]<=16'd4854; ROM2[3895]<=16'd0; ROM3[3895]<=16'd23835; ROM4[3895]<=16'd57324;
ROM1[3896]<=16'd4827; ROM2[3896]<=16'd0; ROM3[3896]<=16'd23826; ROM4[3896]<=16'd57311;
ROM1[3897]<=16'd4823; ROM2[3897]<=16'd0; ROM3[3897]<=16'd23813; ROM4[3897]<=16'd57301;
ROM1[3898]<=16'd4840; ROM2[3898]<=16'd0; ROM3[3898]<=16'd23798; ROM4[3898]<=16'd57295;
ROM1[3899]<=16'd4875; ROM2[3899]<=16'd0; ROM3[3899]<=16'd23792; ROM4[3899]<=16'd57302;
ROM1[3900]<=16'd4889; ROM2[3900]<=16'd0; ROM3[3900]<=16'd23794; ROM4[3900]<=16'd57309;
ROM1[3901]<=16'd4871; ROM2[3901]<=16'd0; ROM3[3901]<=16'd23788; ROM4[3901]<=16'd57299;
ROM1[3902]<=16'd4854; ROM2[3902]<=16'd0; ROM3[3902]<=16'd23783; ROM4[3902]<=16'd57293;
ROM1[3903]<=16'd4849; ROM2[3903]<=16'd0; ROM3[3903]<=16'd23790; ROM4[3903]<=16'd57301;
ROM1[3904]<=16'd4832; ROM2[3904]<=16'd0; ROM3[3904]<=16'd23798; ROM4[3904]<=16'd57309;
ROM1[3905]<=16'd4838; ROM2[3905]<=16'd0; ROM3[3905]<=16'd23808; ROM4[3905]<=16'd57315;
ROM1[3906]<=16'd4885; ROM2[3906]<=16'd0; ROM3[3906]<=16'd23826; ROM4[3906]<=16'd57337;
ROM1[3907]<=16'd4928; ROM2[3907]<=16'd0; ROM3[3907]<=16'd23822; ROM4[3907]<=16'd57344;
ROM1[3908]<=16'd4921; ROM2[3908]<=16'd0; ROM3[3908]<=16'd23798; ROM4[3908]<=16'd57319;
ROM1[3909]<=16'd4909; ROM2[3909]<=16'd0; ROM3[3909]<=16'd23805; ROM4[3909]<=16'd57320;
ROM1[3910]<=16'd4891; ROM2[3910]<=16'd0; ROM3[3910]<=16'd23815; ROM4[3910]<=16'd57325;
ROM1[3911]<=16'd4872; ROM2[3911]<=16'd0; ROM3[3911]<=16'd23812; ROM4[3911]<=16'd57315;
ROM1[3912]<=16'd4868; ROM2[3912]<=16'd0; ROM3[3912]<=16'd23825; ROM4[3912]<=16'd57320;
ROM1[3913]<=16'd4862; ROM2[3913]<=16'd0; ROM3[3913]<=16'd23832; ROM4[3913]<=16'd57326;
ROM1[3914]<=16'd4867; ROM2[3914]<=16'd0; ROM3[3914]<=16'd23823; ROM4[3914]<=16'd57323;
ROM1[3915]<=16'd4891; ROM2[3915]<=16'd0; ROM3[3915]<=16'd23811; ROM4[3915]<=16'd57321;
ROM1[3916]<=16'd4915; ROM2[3916]<=16'd0; ROM3[3916]<=16'd23806; ROM4[3916]<=16'd57323;
ROM1[3917]<=16'd4909; ROM2[3917]<=16'd0; ROM3[3917]<=16'd23808; ROM4[3917]<=16'd57326;
ROM1[3918]<=16'd4890; ROM2[3918]<=16'd0; ROM3[3918]<=16'd23817; ROM4[3918]<=16'd57331;
ROM1[3919]<=16'd4875; ROM2[3919]<=16'd0; ROM3[3919]<=16'd23830; ROM4[3919]<=16'd57334;
ROM1[3920]<=16'd4862; ROM2[3920]<=16'd0; ROM3[3920]<=16'd23836; ROM4[3920]<=16'd57335;
ROM1[3921]<=16'd4858; ROM2[3921]<=16'd0; ROM3[3921]<=16'd23848; ROM4[3921]<=16'd57338;
ROM1[3922]<=16'd4877; ROM2[3922]<=16'd0; ROM3[3922]<=16'd23853; ROM4[3922]<=16'd57341;
ROM1[3923]<=16'd4909; ROM2[3923]<=16'd0; ROM3[3923]<=16'd23849; ROM4[3923]<=16'd57347;
ROM1[3924]<=16'd4943; ROM2[3924]<=16'd0; ROM3[3924]<=16'd23848; ROM4[3924]<=16'd57355;
ROM1[3925]<=16'd4926; ROM2[3925]<=16'd0; ROM3[3925]<=16'd23825; ROM4[3925]<=16'd57337;
ROM1[3926]<=16'd4900; ROM2[3926]<=16'd0; ROM3[3926]<=16'd23825; ROM4[3926]<=16'd57328;
ROM1[3927]<=16'd4891; ROM2[3927]<=16'd0; ROM3[3927]<=16'd23839; ROM4[3927]<=16'd57335;
ROM1[3928]<=16'd4881; ROM2[3928]<=16'd0; ROM3[3928]<=16'd23840; ROM4[3928]<=16'd57337;
ROM1[3929]<=16'd4861; ROM2[3929]<=16'd0; ROM3[3929]<=16'd23840; ROM4[3929]<=16'd57332;
ROM1[3930]<=16'd4854; ROM2[3930]<=16'd0; ROM3[3930]<=16'd23837; ROM4[3930]<=16'd57332;
ROM1[3931]<=16'd4862; ROM2[3931]<=16'd0; ROM3[3931]<=16'd23822; ROM4[3931]<=16'd57328;
ROM1[3932]<=16'd4888; ROM2[3932]<=16'd0; ROM3[3932]<=16'd23802; ROM4[3932]<=16'd57321;
ROM1[3933]<=16'd4911; ROM2[3933]<=16'd0; ROM3[3933]<=16'd23802; ROM4[3933]<=16'd57330;
ROM1[3934]<=16'd4897; ROM2[3934]<=16'd0; ROM3[3934]<=16'd23808; ROM4[3934]<=16'd57331;
ROM1[3935]<=16'd4879; ROM2[3935]<=16'd0; ROM3[3935]<=16'd23815; ROM4[3935]<=16'd57328;
ROM1[3936]<=16'd4866; ROM2[3936]<=16'd0; ROM3[3936]<=16'd23819; ROM4[3936]<=16'd57327;
ROM1[3937]<=16'd4859; ROM2[3937]<=16'd0; ROM3[3937]<=16'd23834; ROM4[3937]<=16'd57332;
ROM1[3938]<=16'd4853; ROM2[3938]<=16'd0; ROM3[3938]<=16'd23839; ROM4[3938]<=16'd57333;
ROM1[3939]<=16'd4855; ROM2[3939]<=16'd0; ROM3[3939]<=16'd23827; ROM4[3939]<=16'd57325;
ROM1[3940]<=16'd4880; ROM2[3940]<=16'd0; ROM3[3940]<=16'd23816; ROM4[3940]<=16'd57321;
ROM1[3941]<=16'd4907; ROM2[3941]<=16'd0; ROM3[3941]<=16'd23813; ROM4[3941]<=16'd57326;
ROM1[3942]<=16'd4912; ROM2[3942]<=16'd0; ROM3[3942]<=16'd23826; ROM4[3942]<=16'd57337;
ROM1[3943]<=16'd4890; ROM2[3943]<=16'd0; ROM3[3943]<=16'd23831; ROM4[3943]<=16'd57332;
ROM1[3944]<=16'd4865; ROM2[3944]<=16'd0; ROM3[3944]<=16'd23833; ROM4[3944]<=16'd57321;
ROM1[3945]<=16'd4850; ROM2[3945]<=16'd0; ROM3[3945]<=16'd23835; ROM4[3945]<=16'd57318;
ROM1[3946]<=16'd4829; ROM2[3946]<=16'd0; ROM3[3946]<=16'd23825; ROM4[3946]<=16'd57307;
ROM1[3947]<=16'd4849; ROM2[3947]<=16'd0; ROM3[3947]<=16'd23834; ROM4[3947]<=16'd57318;
ROM1[3948]<=16'd4891; ROM2[3948]<=16'd0; ROM3[3948]<=16'd23839; ROM4[3948]<=16'd57334;
ROM1[3949]<=16'd4906; ROM2[3949]<=16'd0; ROM3[3949]<=16'd23813; ROM4[3949]<=16'd57323;
ROM1[3950]<=16'd4901; ROM2[3950]<=16'd0; ROM3[3950]<=16'd23804; ROM4[3950]<=16'd57315;
ROM1[3951]<=16'd4877; ROM2[3951]<=16'd0; ROM3[3951]<=16'd23809; ROM4[3951]<=16'd57310;
ROM1[3952]<=16'd4858; ROM2[3952]<=16'd0; ROM3[3952]<=16'd23812; ROM4[3952]<=16'd57309;
ROM1[3953]<=16'd4856; ROM2[3953]<=16'd0; ROM3[3953]<=16'd23826; ROM4[3953]<=16'd57322;
ROM1[3954]<=16'd4850; ROM2[3954]<=16'd0; ROM3[3954]<=16'd23837; ROM4[3954]<=16'd57331;
ROM1[3955]<=16'd4858; ROM2[3955]<=16'd0; ROM3[3955]<=16'd23841; ROM4[3955]<=16'd57337;
ROM1[3956]<=16'd4867; ROM2[3956]<=16'd0; ROM3[3956]<=16'd23824; ROM4[3956]<=16'd57331;
ROM1[3957]<=16'd4882; ROM2[3957]<=16'd0; ROM3[3957]<=16'd23798; ROM4[3957]<=16'd57314;
ROM1[3958]<=16'd4892; ROM2[3958]<=16'd0; ROM3[3958]<=16'd23791; ROM4[3958]<=16'd57314;
ROM1[3959]<=16'd4887; ROM2[3959]<=16'd0; ROM3[3959]<=16'd23797; ROM4[3959]<=16'd57320;
ROM1[3960]<=16'd4886; ROM2[3960]<=16'd0; ROM3[3960]<=16'd23821; ROM4[3960]<=16'd57332;
ROM1[3961]<=16'd4881; ROM2[3961]<=16'd0; ROM3[3961]<=16'd23837; ROM4[3961]<=16'd57341;
ROM1[3962]<=16'd4855; ROM2[3962]<=16'd0; ROM3[3962]<=16'd23830; ROM4[3962]<=16'd57332;
ROM1[3963]<=16'd4838; ROM2[3963]<=16'd0; ROM3[3963]<=16'd23822; ROM4[3963]<=16'd57320;
ROM1[3964]<=16'd4848; ROM2[3964]<=16'd0; ROM3[3964]<=16'd23815; ROM4[3964]<=16'd57319;
ROM1[3965]<=16'd4884; ROM2[3965]<=16'd0; ROM3[3965]<=16'd23805; ROM4[3965]<=16'd57326;
ROM1[3966]<=16'd4906; ROM2[3966]<=16'd0; ROM3[3966]<=16'd23790; ROM4[3966]<=16'd57321;
ROM1[3967]<=16'd4891; ROM2[3967]<=16'd0; ROM3[3967]<=16'd23783; ROM4[3967]<=16'd57312;
ROM1[3968]<=16'd4865; ROM2[3968]<=16'd0; ROM3[3968]<=16'd23789; ROM4[3968]<=16'd57310;
ROM1[3969]<=16'd4860; ROM2[3969]<=16'd0; ROM3[3969]<=16'd23812; ROM4[3969]<=16'd57323;
ROM1[3970]<=16'd4871; ROM2[3970]<=16'd0; ROM3[3970]<=16'd23841; ROM4[3970]<=16'd57347;
ROM1[3971]<=16'd4877; ROM2[3971]<=16'd0; ROM3[3971]<=16'd23859; ROM4[3971]<=16'd57358;
ROM1[3972]<=16'd4883; ROM2[3972]<=16'd0; ROM3[3972]<=16'd23854; ROM4[3972]<=16'd57351;
ROM1[3973]<=16'd4900; ROM2[3973]<=16'd0; ROM3[3973]<=16'd23842; ROM4[3973]<=16'd57343;
ROM1[3974]<=16'd4917; ROM2[3974]<=16'd0; ROM3[3974]<=16'd23831; ROM4[3974]<=16'd57335;
ROM1[3975]<=16'd4912; ROM2[3975]<=16'd0; ROM3[3975]<=16'd23825; ROM4[3975]<=16'd57333;
ROM1[3976]<=16'd4908; ROM2[3976]<=16'd0; ROM3[3976]<=16'd23839; ROM4[3976]<=16'd57346;
ROM1[3977]<=16'd4886; ROM2[3977]<=16'd0; ROM3[3977]<=16'd23842; ROM4[3977]<=16'd57339;
ROM1[3978]<=16'd4865; ROM2[3978]<=16'd0; ROM3[3978]<=16'd23841; ROM4[3978]<=16'd57328;
ROM1[3979]<=16'd4851; ROM2[3979]<=16'd0; ROM3[3979]<=16'd23848; ROM4[3979]<=16'd57327;
ROM1[3980]<=16'd4860; ROM2[3980]<=16'd0; ROM3[3980]<=16'd23854; ROM4[3980]<=16'd57335;
ROM1[3981]<=16'd4901; ROM2[3981]<=16'd0; ROM3[3981]<=16'd23867; ROM4[3981]<=16'd57355;
ROM1[3982]<=16'd4928; ROM2[3982]<=16'd0; ROM3[3982]<=16'd23848; ROM4[3982]<=16'd57349;
ROM1[3983]<=16'd4923; ROM2[3983]<=16'd0; ROM3[3983]<=16'd23821; ROM4[3983]<=16'd57333;
ROM1[3984]<=16'd4909; ROM2[3984]<=16'd0; ROM3[3984]<=16'd23823; ROM4[3984]<=16'd57331;
ROM1[3985]<=16'd4885; ROM2[3985]<=16'd0; ROM3[3985]<=16'd23827; ROM4[3985]<=16'd57326;
ROM1[3986]<=16'd4866; ROM2[3986]<=16'd0; ROM3[3986]<=16'd23827; ROM4[3986]<=16'd57324;
ROM1[3987]<=16'd4848; ROM2[3987]<=16'd0; ROM3[3987]<=16'd23829; ROM4[3987]<=16'd57320;
ROM1[3988]<=16'd4835; ROM2[3988]<=16'd0; ROM3[3988]<=16'd23824; ROM4[3988]<=16'd57315;
ROM1[3989]<=16'd4846; ROM2[3989]<=16'd0; ROM3[3989]<=16'd23812; ROM4[3989]<=16'd57310;
ROM1[3990]<=16'd4884; ROM2[3990]<=16'd0; ROM3[3990]<=16'd23808; ROM4[3990]<=16'd57314;
ROM1[3991]<=16'd4917; ROM2[3991]<=16'd0; ROM3[3991]<=16'd23808; ROM4[3991]<=16'd57327;
ROM1[3992]<=16'd4901; ROM2[3992]<=16'd0; ROM3[3992]<=16'd23803; ROM4[3992]<=16'd57323;
ROM1[3993]<=16'd4883; ROM2[3993]<=16'd0; ROM3[3993]<=16'd23812; ROM4[3993]<=16'd57326;
ROM1[3994]<=16'd4885; ROM2[3994]<=16'd0; ROM3[3994]<=16'd23831; ROM4[3994]<=16'd57341;
ROM1[3995]<=16'd4877; ROM2[3995]<=16'd0; ROM3[3995]<=16'd23844; ROM4[3995]<=16'd57348;
ROM1[3996]<=16'd4864; ROM2[3996]<=16'd0; ROM3[3996]<=16'd23842; ROM4[3996]<=16'd57344;
ROM1[3997]<=16'd4857; ROM2[3997]<=16'd0; ROM3[3997]<=16'd23829; ROM4[3997]<=16'd57326;
ROM1[3998]<=16'd4864; ROM2[3998]<=16'd0; ROM3[3998]<=16'd23802; ROM4[3998]<=16'd57306;
ROM1[3999]<=16'd4889; ROM2[3999]<=16'd0; ROM3[3999]<=16'd23789; ROM4[3999]<=16'd57302;
ROM1[4000]<=16'd4886; ROM2[4000]<=16'd0; ROM3[4000]<=16'd23786; ROM4[4000]<=16'd57295;
ROM1[4001]<=16'd4874; ROM2[4001]<=16'd0; ROM3[4001]<=16'd23791; ROM4[4001]<=16'd57302;
ROM1[4002]<=16'd4863; ROM2[4002]<=16'd0; ROM3[4002]<=16'd23806; ROM4[4002]<=16'd57309;
ROM1[4003]<=16'd4842; ROM2[4003]<=16'd0; ROM3[4003]<=16'd23807; ROM4[4003]<=16'd57304;
ROM1[4004]<=16'd4824; ROM2[4004]<=16'd0; ROM3[4004]<=16'd23810; ROM4[4004]<=16'd57305;
ROM1[4005]<=16'd4829; ROM2[4005]<=16'd0; ROM3[4005]<=16'd23818; ROM4[4005]<=16'd57310;
ROM1[4006]<=16'd4858; ROM2[4006]<=16'd0; ROM3[4006]<=16'd23818; ROM4[4006]<=16'd57318;
ROM1[4007]<=16'd4891; ROM2[4007]<=16'd0; ROM3[4007]<=16'd23804; ROM4[4007]<=16'd57319;
ROM1[4008]<=16'd4904; ROM2[4008]<=16'd0; ROM3[4008]<=16'd23799; ROM4[4008]<=16'd57319;
ROM1[4009]<=16'd4890; ROM2[4009]<=16'd0; ROM3[4009]<=16'd23801; ROM4[4009]<=16'd57317;
ROM1[4010]<=16'd4863; ROM2[4010]<=16'd0; ROM3[4010]<=16'd23800; ROM4[4010]<=16'd57312;
ROM1[4011]<=16'd4849; ROM2[4011]<=16'd0; ROM3[4011]<=16'd23811; ROM4[4011]<=16'd57314;
ROM1[4012]<=16'd4844; ROM2[4012]<=16'd0; ROM3[4012]<=16'd23822; ROM4[4012]<=16'd57315;
ROM1[4013]<=16'd4837; ROM2[4013]<=16'd0; ROM3[4013]<=16'd23820; ROM4[4013]<=16'd57312;
ROM1[4014]<=16'd4859; ROM2[4014]<=16'd0; ROM3[4014]<=16'd23828; ROM4[4014]<=16'd57321;
ROM1[4015]<=16'd4913; ROM2[4015]<=16'd0; ROM3[4015]<=16'd23843; ROM4[4015]<=16'd57349;
ROM1[4016]<=16'd4932; ROM2[4016]<=16'd0; ROM3[4016]<=16'd23832; ROM4[4016]<=16'd57350;
ROM1[4017]<=16'd4905; ROM2[4017]<=16'd0; ROM3[4017]<=16'd23815; ROM4[4017]<=16'd57332;
ROM1[4018]<=16'd4869; ROM2[4018]<=16'd0; ROM3[4018]<=16'd23807; ROM4[4018]<=16'd57319;
ROM1[4019]<=16'd4844; ROM2[4019]<=16'd0; ROM3[4019]<=16'd23807; ROM4[4019]<=16'd57310;
ROM1[4020]<=16'd4837; ROM2[4020]<=16'd0; ROM3[4020]<=16'd23813; ROM4[4020]<=16'd57310;
ROM1[4021]<=16'd4830; ROM2[4021]<=16'd0; ROM3[4021]<=16'd23818; ROM4[4021]<=16'd57311;
ROM1[4022]<=16'd4838; ROM2[4022]<=16'd0; ROM3[4022]<=16'd23818; ROM4[4022]<=16'd57308;
ROM1[4023]<=16'd4865; ROM2[4023]<=16'd0; ROM3[4023]<=16'd23808; ROM4[4023]<=16'd57307;
ROM1[4024]<=16'd4886; ROM2[4024]<=16'd0; ROM3[4024]<=16'd23789; ROM4[4024]<=16'd57301;
ROM1[4025]<=16'd4887; ROM2[4025]<=16'd0; ROM3[4025]<=16'd23787; ROM4[4025]<=16'd57298;
ROM1[4026]<=16'd4878; ROM2[4026]<=16'd0; ROM3[4026]<=16'd23793; ROM4[4026]<=16'd57305;
ROM1[4027]<=16'd4868; ROM2[4027]<=16'd0; ROM3[4027]<=16'd23812; ROM4[4027]<=16'd57314;
ROM1[4028]<=16'd4854; ROM2[4028]<=16'd0; ROM3[4028]<=16'd23820; ROM4[4028]<=16'd57315;
ROM1[4029]<=16'd4826; ROM2[4029]<=16'd0; ROM3[4029]<=16'd23812; ROM4[4029]<=16'd57304;
ROM1[4030]<=16'd4827; ROM2[4030]<=16'd0; ROM3[4030]<=16'd23808; ROM4[4030]<=16'd57304;
ROM1[4031]<=16'd4849; ROM2[4031]<=16'd0; ROM3[4031]<=16'd23791; ROM4[4031]<=16'd57299;
ROM1[4032]<=16'd4898; ROM2[4032]<=16'd0; ROM3[4032]<=16'd23799; ROM4[4032]<=16'd57312;
ROM1[4033]<=16'd4911; ROM2[4033]<=16'd0; ROM3[4033]<=16'd23801; ROM4[4033]<=16'd57318;
ROM1[4034]<=16'd4866; ROM2[4034]<=16'd0; ROM3[4034]<=16'd23785; ROM4[4034]<=16'd57293;
ROM1[4035]<=16'd4836; ROM2[4035]<=16'd0; ROM3[4035]<=16'd23788; ROM4[4035]<=16'd57284;
ROM1[4036]<=16'd4818; ROM2[4036]<=16'd0; ROM3[4036]<=16'd23791; ROM4[4036]<=16'd57283;
ROM1[4037]<=16'd4813; ROM2[4037]<=16'd0; ROM3[4037]<=16'd23807; ROM4[4037]<=16'd57292;
ROM1[4038]<=16'd4827; ROM2[4038]<=16'd0; ROM3[4038]<=16'd23830; ROM4[4038]<=16'd57309;
ROM1[4039]<=16'd4834; ROM2[4039]<=16'd0; ROM3[4039]<=16'd23820; ROM4[4039]<=16'd57302;
ROM1[4040]<=16'd4854; ROM2[4040]<=16'd0; ROM3[4040]<=16'd23796; ROM4[4040]<=16'd57289;
ROM1[4041]<=16'd4885; ROM2[4041]<=16'd0; ROM3[4041]<=16'd23790; ROM4[4041]<=16'd57294;
ROM1[4042]<=16'd4888; ROM2[4042]<=16'd0; ROM3[4042]<=16'd23795; ROM4[4042]<=16'd57297;
ROM1[4043]<=16'd4873; ROM2[4043]<=16'd0; ROM3[4043]<=16'd23806; ROM4[4043]<=16'd57301;
ROM1[4044]<=16'd4862; ROM2[4044]<=16'd0; ROM3[4044]<=16'd23821; ROM4[4044]<=16'd57305;
ROM1[4045]<=16'd4851; ROM2[4045]<=16'd0; ROM3[4045]<=16'd23831; ROM4[4045]<=16'd57307;
ROM1[4046]<=16'd4837; ROM2[4046]<=16'd0; ROM3[4046]<=16'd23833; ROM4[4046]<=16'd57306;
ROM1[4047]<=16'd4848; ROM2[4047]<=16'd0; ROM3[4047]<=16'd23834; ROM4[4047]<=16'd57313;
ROM1[4048]<=16'd4870; ROM2[4048]<=16'd0; ROM3[4048]<=16'd23818; ROM4[4048]<=16'd57309;
ROM1[4049]<=16'd4890; ROM2[4049]<=16'd0; ROM3[4049]<=16'd23794; ROM4[4049]<=16'd57304;
ROM1[4050]<=16'd4902; ROM2[4050]<=16'd0; ROM3[4050]<=16'd23801; ROM4[4050]<=16'd57315;
ROM1[4051]<=16'd4888; ROM2[4051]<=16'd0; ROM3[4051]<=16'd23806; ROM4[4051]<=16'd57314;
ROM1[4052]<=16'd4862; ROM2[4052]<=16'd0; ROM3[4052]<=16'd23801; ROM4[4052]<=16'd57309;
ROM1[4053]<=16'd4853; ROM2[4053]<=16'd0; ROM3[4053]<=16'd23809; ROM4[4053]<=16'd57310;
ROM1[4054]<=16'd4843; ROM2[4054]<=16'd0; ROM3[4054]<=16'd23820; ROM4[4054]<=16'd57311;
ROM1[4055]<=16'd4835; ROM2[4055]<=16'd0; ROM3[4055]<=16'd23811; ROM4[4055]<=16'd57304;
ROM1[4056]<=16'd4858; ROM2[4056]<=16'd0; ROM3[4056]<=16'd23806; ROM4[4056]<=16'd57307;
ROM1[4057]<=16'd4892; ROM2[4057]<=16'd0; ROM3[4057]<=16'd23800; ROM4[4057]<=16'd57313;
ROM1[4058]<=16'd4894; ROM2[4058]<=16'd0; ROM3[4058]<=16'd23790; ROM4[4058]<=16'd57304;
ROM1[4059]<=16'd4878; ROM2[4059]<=16'd0; ROM3[4059]<=16'd23797; ROM4[4059]<=16'd57304;
ROM1[4060]<=16'd4861; ROM2[4060]<=16'd0; ROM3[4060]<=16'd23809; ROM4[4060]<=16'd57308;
ROM1[4061]<=16'd4847; ROM2[4061]<=16'd0; ROM3[4061]<=16'd23815; ROM4[4061]<=16'd57307;
ROM1[4062]<=16'd4827; ROM2[4062]<=16'd0; ROM3[4062]<=16'd23811; ROM4[4062]<=16'd57300;
ROM1[4063]<=16'd4816; ROM2[4063]<=16'd0; ROM3[4063]<=16'd23806; ROM4[4063]<=16'd57291;
ROM1[4064]<=16'd4825; ROM2[4064]<=16'd0; ROM3[4064]<=16'd23801; ROM4[4064]<=16'd57288;
ROM1[4065]<=16'd4854; ROM2[4065]<=16'd0; ROM3[4065]<=16'd23787; ROM4[4065]<=16'd57286;
ROM1[4066]<=16'd4887; ROM2[4066]<=16'd0; ROM3[4066]<=16'd23781; ROM4[4066]<=16'd57295;
ROM1[4067]<=16'd4873; ROM2[4067]<=16'd0; ROM3[4067]<=16'd23776; ROM4[4067]<=16'd57292;
ROM1[4068]<=16'd4847; ROM2[4068]<=16'd0; ROM3[4068]<=16'd23775; ROM4[4068]<=16'd57286;
ROM1[4069]<=16'd4839; ROM2[4069]<=16'd0; ROM3[4069]<=16'd23788; ROM4[4069]<=16'd57290;
ROM1[4070]<=16'd4831; ROM2[4070]<=16'd0; ROM3[4070]<=16'd23804; ROM4[4070]<=16'd57296;
ROM1[4071]<=16'd4824; ROM2[4071]<=16'd0; ROM3[4071]<=16'd23812; ROM4[4071]<=16'd57298;
ROM1[4072]<=16'd4839; ROM2[4072]<=16'd0; ROM3[4072]<=16'd23816; ROM4[4072]<=16'd57302;
ROM1[4073]<=16'd4868; ROM2[4073]<=16'd0; ROM3[4073]<=16'd23808; ROM4[4073]<=16'd57303;
ROM1[4074]<=16'd4894; ROM2[4074]<=16'd0; ROM3[4074]<=16'd23793; ROM4[4074]<=16'd57302;
ROM1[4075]<=16'd4903; ROM2[4075]<=16'd0; ROM3[4075]<=16'd23795; ROM4[4075]<=16'd57310;
ROM1[4076]<=16'd4884; ROM2[4076]<=16'd0; ROM3[4076]<=16'd23798; ROM4[4076]<=16'd57312;
ROM1[4077]<=16'd4855; ROM2[4077]<=16'd0; ROM3[4077]<=16'd23798; ROM4[4077]<=16'd57309;
ROM1[4078]<=16'd4836; ROM2[4078]<=16'd0; ROM3[4078]<=16'd23796; ROM4[4078]<=16'd57304;
ROM1[4079]<=16'd4822; ROM2[4079]<=16'd0; ROM3[4079]<=16'd23798; ROM4[4079]<=16'd57300;
ROM1[4080]<=16'd4840; ROM2[4080]<=16'd0; ROM3[4080]<=16'd23809; ROM4[4080]<=16'd57313;
ROM1[4081]<=16'd4862; ROM2[4081]<=16'd0; ROM3[4081]<=16'd23804; ROM4[4081]<=16'd57313;
ROM1[4082]<=16'd4877; ROM2[4082]<=16'd0; ROM3[4082]<=16'd23773; ROM4[4082]<=16'd57296;
ROM1[4083]<=16'd4883; ROM2[4083]<=16'd0; ROM3[4083]<=16'd23760; ROM4[4083]<=16'd57289;
ROM1[4084]<=16'd4867; ROM2[4084]<=16'd0; ROM3[4084]<=16'd23771; ROM4[4084]<=16'd57294;
ROM1[4085]<=16'd4874; ROM2[4085]<=16'd0; ROM3[4085]<=16'd23804; ROM4[4085]<=16'd57319;
ROM1[4086]<=16'd4869; ROM2[4086]<=16'd0; ROM3[4086]<=16'd23821; ROM4[4086]<=16'd57328;
ROM1[4087]<=16'd4839; ROM2[4087]<=16'd0; ROM3[4087]<=16'd23816; ROM4[4087]<=16'd57315;
ROM1[4088]<=16'd4834; ROM2[4088]<=16'd0; ROM3[4088]<=16'd23814; ROM4[4088]<=16'd57310;
ROM1[4089]<=16'd4838; ROM2[4089]<=16'd0; ROM3[4089]<=16'd23805; ROM4[4089]<=16'd57300;
ROM1[4090]<=16'd4864; ROM2[4090]<=16'd0; ROM3[4090]<=16'd23801; ROM4[4090]<=16'd57301;
ROM1[4091]<=16'd4898; ROM2[4091]<=16'd0; ROM3[4091]<=16'd23805; ROM4[4091]<=16'd57316;
ROM1[4092]<=16'd4896; ROM2[4092]<=16'd0; ROM3[4092]<=16'd23809; ROM4[4092]<=16'd57318;
ROM1[4093]<=16'd4869; ROM2[4093]<=16'd0; ROM3[4093]<=16'd23806; ROM4[4093]<=16'd57309;
ROM1[4094]<=16'd4865; ROM2[4094]<=16'd0; ROM3[4094]<=16'd23829; ROM4[4094]<=16'd57321;
ROM1[4095]<=16'd4854; ROM2[4095]<=16'd0; ROM3[4095]<=16'd23844; ROM4[4095]<=16'd57327;
ROM1[4096]<=16'd4820; ROM2[4096]<=16'd0; ROM3[4096]<=16'd23831; ROM4[4096]<=16'd57310;
ROM1[4097]<=16'd4827; ROM2[4097]<=16'd0; ROM3[4097]<=16'd23828; ROM4[4097]<=16'd57310;
ROM1[4098]<=16'd4863; ROM2[4098]<=16'd0; ROM3[4098]<=16'd23819; ROM4[4098]<=16'd57313;
ROM1[4099]<=16'd4910; ROM2[4099]<=16'd0; ROM3[4099]<=16'd23826; ROM4[4099]<=16'd57331;
ROM1[4100]<=16'd4907; ROM2[4100]<=16'd0; ROM3[4100]<=16'd23821; ROM4[4100]<=16'd57328;
ROM1[4101]<=16'd4873; ROM2[4101]<=16'd0; ROM3[4101]<=16'd23815; ROM4[4101]<=16'd57310;
ROM1[4102]<=16'd4861; ROM2[4102]<=16'd0; ROM3[4102]<=16'd23829; ROM4[4102]<=16'd57317;
ROM1[4103]<=16'd4850; ROM2[4103]<=16'd0; ROM3[4103]<=16'd23833; ROM4[4103]<=16'd57317;
ROM1[4104]<=16'd4845; ROM2[4104]<=16'd0; ROM3[4104]<=16'd23842; ROM4[4104]<=16'd57323;
ROM1[4105]<=16'd4856; ROM2[4105]<=16'd0; ROM3[4105]<=16'd23852; ROM4[4105]<=16'd57335;
ROM1[4106]<=16'd4874; ROM2[4106]<=16'd0; ROM3[4106]<=16'd23848; ROM4[4106]<=16'd57335;
ROM1[4107]<=16'd4898; ROM2[4107]<=16'd0; ROM3[4107]<=16'd23833; ROM4[4107]<=16'd57334;
ROM1[4108]<=16'd4924; ROM2[4108]<=16'd0; ROM3[4108]<=16'd23843; ROM4[4108]<=16'd57349;
ROM1[4109]<=16'd4925; ROM2[4109]<=16'd0; ROM3[4109]<=16'd23856; ROM4[4109]<=16'd57362;
ROM1[4110]<=16'd4898; ROM2[4110]<=16'd0; ROM3[4110]<=16'd23849; ROM4[4110]<=16'd57351;
ROM1[4111]<=16'd4880; ROM2[4111]<=16'd0; ROM3[4111]<=16'd23843; ROM4[4111]<=16'd57340;
ROM1[4112]<=16'd4862; ROM2[4112]<=16'd0; ROM3[4112]<=16'd23844; ROM4[4112]<=16'd57337;
ROM1[4113]<=16'd4841; ROM2[4113]<=16'd0; ROM3[4113]<=16'd23836; ROM4[4113]<=16'd57323;
ROM1[4114]<=16'd4851; ROM2[4114]<=16'd0; ROM3[4114]<=16'd23830; ROM4[4114]<=16'd57318;
ROM1[4115]<=16'd4883; ROM2[4115]<=16'd0; ROM3[4115]<=16'd23824; ROM4[4115]<=16'd57322;
ROM1[4116]<=16'd4900; ROM2[4116]<=16'd0; ROM3[4116]<=16'd23813; ROM4[4116]<=16'd57318;
ROM1[4117]<=16'd4891; ROM2[4117]<=16'd0; ROM3[4117]<=16'd23814; ROM4[4117]<=16'd57318;
ROM1[4118]<=16'd4872; ROM2[4118]<=16'd0; ROM3[4118]<=16'd23815; ROM4[4118]<=16'd57317;
ROM1[4119]<=16'd4854; ROM2[4119]<=16'd0; ROM3[4119]<=16'd23818; ROM4[4119]<=16'd57313;
ROM1[4120]<=16'd4834; ROM2[4120]<=16'd0; ROM3[4120]<=16'd23820; ROM4[4120]<=16'd57309;
ROM1[4121]<=16'd4835; ROM2[4121]<=16'd0; ROM3[4121]<=16'd23831; ROM4[4121]<=16'd57320;
ROM1[4122]<=16'd4850; ROM2[4122]<=16'd0; ROM3[4122]<=16'd23835; ROM4[4122]<=16'd57328;
ROM1[4123]<=16'd4873; ROM2[4123]<=16'd0; ROM3[4123]<=16'd23822; ROM4[4123]<=16'd57323;
ROM1[4124]<=16'd4904; ROM2[4124]<=16'd0; ROM3[4124]<=16'd23811; ROM4[4124]<=16'd57321;
ROM1[4125]<=16'd4895; ROM2[4125]<=16'd0; ROM3[4125]<=16'd23804; ROM4[4125]<=16'd57316;
ROM1[4126]<=16'd4874; ROM2[4126]<=16'd0; ROM3[4126]<=16'd23808; ROM4[4126]<=16'd57317;
ROM1[4127]<=16'd4869; ROM2[4127]<=16'd0; ROM3[4127]<=16'd23828; ROM4[4127]<=16'd57328;
ROM1[4128]<=16'd4859; ROM2[4128]<=16'd0; ROM3[4128]<=16'd23834; ROM4[4128]<=16'd57329;
ROM1[4129]<=16'd4845; ROM2[4129]<=16'd0; ROM3[4129]<=16'd23837; ROM4[4129]<=16'd57327;
ROM1[4130]<=16'd4848; ROM2[4130]<=16'd0; ROM3[4130]<=16'd23840; ROM4[4130]<=16'd57328;
ROM1[4131]<=16'd4879; ROM2[4131]<=16'd0; ROM3[4131]<=16'd23843; ROM4[4131]<=16'd57342;
ROM1[4132]<=16'd4914; ROM2[4132]<=16'd0; ROM3[4132]<=16'd23832; ROM4[4132]<=16'd57339;
ROM1[4133]<=16'd4902; ROM2[4133]<=16'd0; ROM3[4133]<=16'd23803; ROM4[4133]<=16'd57311;
ROM1[4134]<=16'd4880; ROM2[4134]<=16'd0; ROM3[4134]<=16'd23804; ROM4[4134]<=16'd57308;
ROM1[4135]<=16'd4854; ROM2[4135]<=16'd0; ROM3[4135]<=16'd23807; ROM4[4135]<=16'd57301;
ROM1[4136]<=16'd4842; ROM2[4136]<=16'd0; ROM3[4136]<=16'd23817; ROM4[4136]<=16'd57302;
ROM1[4137]<=16'd4842; ROM2[4137]<=16'd0; ROM3[4137]<=16'd23838; ROM4[4137]<=16'd57318;
ROM1[4138]<=16'd4832; ROM2[4138]<=16'd0; ROM3[4138]<=16'd23831; ROM4[4138]<=16'd57311;
ROM1[4139]<=16'd4832; ROM2[4139]<=16'd0; ROM3[4139]<=16'd23807; ROM4[4139]<=16'd57291;
ROM1[4140]<=16'd4855; ROM2[4140]<=16'd0; ROM3[4140]<=16'd23786; ROM4[4140]<=16'd57284;
ROM1[4141]<=16'd4880; ROM2[4141]<=16'd0; ROM3[4141]<=16'd23780; ROM4[4141]<=16'd57292;
ROM1[4142]<=16'd4899; ROM2[4142]<=16'd0; ROM3[4142]<=16'd23799; ROM4[4142]<=16'd57312;
ROM1[4143]<=16'd4887; ROM2[4143]<=16'd0; ROM3[4143]<=16'd23808; ROM4[4143]<=16'd57319;
ROM1[4144]<=16'd4858; ROM2[4144]<=16'd0; ROM3[4144]<=16'd23808; ROM4[4144]<=16'd57311;
ROM1[4145]<=16'd4842; ROM2[4145]<=16'd0; ROM3[4145]<=16'd23813; ROM4[4145]<=16'd57308;
ROM1[4146]<=16'd4823; ROM2[4146]<=16'd0; ROM3[4146]<=16'd23809; ROM4[4146]<=16'd57300;
ROM1[4147]<=16'd4820; ROM2[4147]<=16'd0; ROM3[4147]<=16'd23803; ROM4[4147]<=16'd57294;
ROM1[4148]<=16'd4846; ROM2[4148]<=16'd0; ROM3[4148]<=16'd23790; ROM4[4148]<=16'd57290;
ROM1[4149]<=16'd4876; ROM2[4149]<=16'd0; ROM3[4149]<=16'd23777; ROM4[4149]<=16'd57289;
ROM1[4150]<=16'd4873; ROM2[4150]<=16'd0; ROM3[4150]<=16'd23775; ROM4[4150]<=16'd57284;
ROM1[4151]<=16'd4860; ROM2[4151]<=16'd0; ROM3[4151]<=16'd23788; ROM4[4151]<=16'd57286;
ROM1[4152]<=16'd4847; ROM2[4152]<=16'd0; ROM3[4152]<=16'd23803; ROM4[4152]<=16'd57295;
ROM1[4153]<=16'd4837; ROM2[4153]<=16'd0; ROM3[4153]<=16'd23811; ROM4[4153]<=16'd57296;
ROM1[4154]<=16'd4826; ROM2[4154]<=16'd0; ROM3[4154]<=16'd23813; ROM4[4154]<=16'd57292;
ROM1[4155]<=16'd4828; ROM2[4155]<=16'd0; ROM3[4155]<=16'd23813; ROM4[4155]<=16'd57297;
ROM1[4156]<=16'd4856; ROM2[4156]<=16'd0; ROM3[4156]<=16'd23814; ROM4[4156]<=16'd57304;
ROM1[4157]<=16'd4888; ROM2[4157]<=16'd0; ROM3[4157]<=16'd23802; ROM4[4157]<=16'd57303;
ROM1[4158]<=16'd4888; ROM2[4158]<=16'd0; ROM3[4158]<=16'd23794; ROM4[4158]<=16'd57296;
ROM1[4159]<=16'd4874; ROM2[4159]<=16'd0; ROM3[4159]<=16'd23796; ROM4[4159]<=16'd57292;
ROM1[4160]<=16'd4863; ROM2[4160]<=16'd0; ROM3[4160]<=16'd23810; ROM4[4160]<=16'd57302;
ROM1[4161]<=16'd4849; ROM2[4161]<=16'd0; ROM3[4161]<=16'd23819; ROM4[4161]<=16'd57303;
ROM1[4162]<=16'd4822; ROM2[4162]<=16'd0; ROM3[4162]<=16'd23814; ROM4[4162]<=16'd57290;
ROM1[4163]<=16'd4807; ROM2[4163]<=16'd0; ROM3[4163]<=16'd23803; ROM4[4163]<=16'd57279;
ROM1[4164]<=16'd4815; ROM2[4164]<=16'd0; ROM3[4164]<=16'd23791; ROM4[4164]<=16'd57271;
ROM1[4165]<=16'd4853; ROM2[4165]<=16'd0; ROM3[4165]<=16'd23785; ROM4[4165]<=16'd57277;
ROM1[4166]<=16'd4880; ROM2[4166]<=16'd0; ROM3[4166]<=16'd23781; ROM4[4166]<=16'd57287;
ROM1[4167]<=16'd4869; ROM2[4167]<=16'd0; ROM3[4167]<=16'd23782; ROM4[4167]<=16'd57285;
ROM1[4168]<=16'd4843; ROM2[4168]<=16'd0; ROM3[4168]<=16'd23780; ROM4[4168]<=16'd57279;
ROM1[4169]<=16'd4822; ROM2[4169]<=16'd0; ROM3[4169]<=16'd23782; ROM4[4169]<=16'd57276;
ROM1[4170]<=16'd4815; ROM2[4170]<=16'd0; ROM3[4170]<=16'd23794; ROM4[4170]<=16'd57280;
ROM1[4171]<=16'd4810; ROM2[4171]<=16'd0; ROM3[4171]<=16'd23799; ROM4[4171]<=16'd57281;
ROM1[4172]<=16'd4819; ROM2[4172]<=16'd0; ROM3[4172]<=16'd23797; ROM4[4172]<=16'd57282;
ROM1[4173]<=16'd4846; ROM2[4173]<=16'd0; ROM3[4173]<=16'd23787; ROM4[4173]<=16'd57281;
ROM1[4174]<=16'd4875; ROM2[4174]<=16'd0; ROM3[4174]<=16'd23777; ROM4[4174]<=16'd57281;
ROM1[4175]<=16'd4881; ROM2[4175]<=16'd0; ROM3[4175]<=16'd23784; ROM4[4175]<=16'd57294;
ROM1[4176]<=16'd4866; ROM2[4176]<=16'd0; ROM3[4176]<=16'd23794; ROM4[4176]<=16'd57299;
ROM1[4177]<=16'd4853; ROM2[4177]<=16'd0; ROM3[4177]<=16'd23805; ROM4[4177]<=16'd57301;
ROM1[4178]<=16'd4847; ROM2[4178]<=16'd0; ROM3[4178]<=16'd23812; ROM4[4178]<=16'd57306;
ROM1[4179]<=16'd4840; ROM2[4179]<=16'd0; ROM3[4179]<=16'd23832; ROM4[4179]<=16'd57315;
ROM1[4180]<=16'd4859; ROM2[4180]<=16'd0; ROM3[4180]<=16'd23853; ROM4[4180]<=16'd57334;
ROM1[4181]<=16'd4880; ROM2[4181]<=16'd0; ROM3[4181]<=16'd23848; ROM4[4181]<=16'd57338;
ROM1[4182]<=16'd4891; ROM2[4182]<=16'd0; ROM3[4182]<=16'd23820; ROM4[4182]<=16'd57322;
ROM1[4183]<=16'd4887; ROM2[4183]<=16'd0; ROM3[4183]<=16'd23801; ROM4[4183]<=16'd57308;
ROM1[4184]<=16'd4865; ROM2[4184]<=16'd0; ROM3[4184]<=16'd23804; ROM4[4184]<=16'd57302;
ROM1[4185]<=16'd4853; ROM2[4185]<=16'd0; ROM3[4185]<=16'd23814; ROM4[4185]<=16'd57307;
ROM1[4186]<=16'd4862; ROM2[4186]<=16'd0; ROM3[4186]<=16'd23841; ROM4[4186]<=16'd57329;
ROM1[4187]<=16'd4851; ROM2[4187]<=16'd0; ROM3[4187]<=16'd23854; ROM4[4187]<=16'd57334;
ROM1[4188]<=16'd4841; ROM2[4188]<=16'd0; ROM3[4188]<=16'd23850; ROM4[4188]<=16'd57327;
ROM1[4189]<=16'd4851; ROM2[4189]<=16'd0; ROM3[4189]<=16'd23837; ROM4[4189]<=16'd57321;
ROM1[4190]<=16'd4877; ROM2[4190]<=16'd0; ROM3[4190]<=16'd23817; ROM4[4190]<=16'd57311;
ROM1[4191]<=16'd4899; ROM2[4191]<=16'd0; ROM3[4191]<=16'd23801; ROM4[4191]<=16'd57307;
ROM1[4192]<=16'd4884; ROM2[4192]<=16'd0; ROM3[4192]<=16'd23789; ROM4[4192]<=16'd57299;
ROM1[4193]<=16'd4859; ROM2[4193]<=16'd0; ROM3[4193]<=16'd23793; ROM4[4193]<=16'd57297;
ROM1[4194]<=16'd4842; ROM2[4194]<=16'd0; ROM3[4194]<=16'd23804; ROM4[4194]<=16'd57302;
ROM1[4195]<=16'd4825; ROM2[4195]<=16'd0; ROM3[4195]<=16'd23804; ROM4[4195]<=16'd57300;
ROM1[4196]<=16'd4823; ROM2[4196]<=16'd0; ROM3[4196]<=16'd23806; ROM4[4196]<=16'd57300;
ROM1[4197]<=16'd4832; ROM2[4197]<=16'd0; ROM3[4197]<=16'd23809; ROM4[4197]<=16'd57304;
ROM1[4198]<=16'd4850; ROM2[4198]<=16'd0; ROM3[4198]<=16'd23798; ROM4[4198]<=16'd57300;
ROM1[4199]<=16'd4881; ROM2[4199]<=16'd0; ROM3[4199]<=16'd23788; ROM4[4199]<=16'd57304;
ROM1[4200]<=16'd4890; ROM2[4200]<=16'd0; ROM3[4200]<=16'd23796; ROM4[4200]<=16'd57310;
ROM1[4201]<=16'd4877; ROM2[4201]<=16'd0; ROM3[4201]<=16'd23804; ROM4[4201]<=16'd57314;
ROM1[4202]<=16'd4862; ROM2[4202]<=16'd0; ROM3[4202]<=16'd23818; ROM4[4202]<=16'd57319;
ROM1[4203]<=16'd4845; ROM2[4203]<=16'd0; ROM3[4203]<=16'd23821; ROM4[4203]<=16'd57315;
ROM1[4204]<=16'd4828; ROM2[4204]<=16'd0; ROM3[4204]<=16'd23820; ROM4[4204]<=16'd57310;
ROM1[4205]<=16'd4828; ROM2[4205]<=16'd0; ROM3[4205]<=16'd23818; ROM4[4205]<=16'd57303;
ROM1[4206]<=16'd4849; ROM2[4206]<=16'd0; ROM3[4206]<=16'd23807; ROM4[4206]<=16'd57300;
ROM1[4207]<=16'd4889; ROM2[4207]<=16'd0; ROM3[4207]<=16'd23806; ROM4[4207]<=16'd57315;
ROM1[4208]<=16'd4897; ROM2[4208]<=16'd0; ROM3[4208]<=16'd23802; ROM4[4208]<=16'd57316;
ROM1[4209]<=16'd4875; ROM2[4209]<=16'd0; ROM3[4209]<=16'd23797; ROM4[4209]<=16'd57307;
ROM1[4210]<=16'd4860; ROM2[4210]<=16'd0; ROM3[4210]<=16'd23802; ROM4[4210]<=16'd57308;
ROM1[4211]<=16'd4849; ROM2[4211]<=16'd0; ROM3[4211]<=16'd23807; ROM4[4211]<=16'd57302;
ROM1[4212]<=16'd4834; ROM2[4212]<=16'd0; ROM3[4212]<=16'd23812; ROM4[4212]<=16'd57303;
ROM1[4213]<=16'd4842; ROM2[4213]<=16'd0; ROM3[4213]<=16'd23828; ROM4[4213]<=16'd57323;
ROM1[4214]<=16'd4863; ROM2[4214]<=16'd0; ROM3[4214]<=16'd23832; ROM4[4214]<=16'd57332;
ROM1[4215]<=16'd4892; ROM2[4215]<=16'd0; ROM3[4215]<=16'd23818; ROM4[4215]<=16'd57329;
ROM1[4216]<=16'd4915; ROM2[4216]<=16'd0; ROM3[4216]<=16'd23808; ROM4[4216]<=16'd57327;
ROM1[4217]<=16'd4891; ROM2[4217]<=16'd0; ROM3[4217]<=16'd23798; ROM4[4217]<=16'd57314;
ROM1[4218]<=16'd4858; ROM2[4218]<=16'd0; ROM3[4218]<=16'd23788; ROM4[4218]<=16'd57301;
ROM1[4219]<=16'd4845; ROM2[4219]<=16'd0; ROM3[4219]<=16'd23793; ROM4[4219]<=16'd57302;
ROM1[4220]<=16'd4829; ROM2[4220]<=16'd0; ROM3[4220]<=16'd23801; ROM4[4220]<=16'd57302;
ROM1[4221]<=16'd4821; ROM2[4221]<=16'd0; ROM3[4221]<=16'd23808; ROM4[4221]<=16'd57304;
ROM1[4222]<=16'd4832; ROM2[4222]<=16'd0; ROM3[4222]<=16'd23810; ROM4[4222]<=16'd57306;
ROM1[4223]<=16'd4870; ROM2[4223]<=16'd0; ROM3[4223]<=16'd23818; ROM4[4223]<=16'd57323;
ROM1[4224]<=16'd4897; ROM2[4224]<=16'd0; ROM3[4224]<=16'd23807; ROM4[4224]<=16'd57322;
ROM1[4225]<=16'd4877; ROM2[4225]<=16'd0; ROM3[4225]<=16'd23785; ROM4[4225]<=16'd57303;
ROM1[4226]<=16'd4856; ROM2[4226]<=16'd0; ROM3[4226]<=16'd23792; ROM4[4226]<=16'd57301;
ROM1[4227]<=16'd4839; ROM2[4227]<=16'd0; ROM3[4227]<=16'd23802; ROM4[4227]<=16'd57303;
ROM1[4228]<=16'd4834; ROM2[4228]<=16'd0; ROM3[4228]<=16'd23812; ROM4[4228]<=16'd57314;
ROM1[4229]<=16'd4817; ROM2[4229]<=16'd0; ROM3[4229]<=16'd23813; ROM4[4229]<=16'd57308;
ROM1[4230]<=16'd4828; ROM2[4230]<=16'd0; ROM3[4230]<=16'd23826; ROM4[4230]<=16'd57316;
ROM1[4231]<=16'd4864; ROM2[4231]<=16'd0; ROM3[4231]<=16'd23843; ROM4[4231]<=16'd57333;
ROM1[4232]<=16'd4879; ROM2[4232]<=16'd0; ROM3[4232]<=16'd23816; ROM4[4232]<=16'd57320;
ROM1[4233]<=16'd4886; ROM2[4233]<=16'd0; ROM3[4233]<=16'd23803; ROM4[4233]<=16'd57312;
ROM1[4234]<=16'd4867; ROM2[4234]<=16'd0; ROM3[4234]<=16'd23796; ROM4[4234]<=16'd57304;
ROM1[4235]<=16'd4834; ROM2[4235]<=16'd0; ROM3[4235]<=16'd23783; ROM4[4235]<=16'd57287;
ROM1[4236]<=16'd4826; ROM2[4236]<=16'd0; ROM3[4236]<=16'd23794; ROM4[4236]<=16'd57291;
ROM1[4237]<=16'd4824; ROM2[4237]<=16'd0; ROM3[4237]<=16'd23813; ROM4[4237]<=16'd57301;
ROM1[4238]<=16'd4832; ROM2[4238]<=16'd0; ROM3[4238]<=16'd23821; ROM4[4238]<=16'd57310;
ROM1[4239]<=16'd4848; ROM2[4239]<=16'd0; ROM3[4239]<=16'd23809; ROM4[4239]<=16'd57309;
ROM1[4240]<=16'd4876; ROM2[4240]<=16'd0; ROM3[4240]<=16'd23800; ROM4[4240]<=16'd57308;
ROM1[4241]<=16'd4902; ROM2[4241]<=16'd0; ROM3[4241]<=16'd23801; ROM4[4241]<=16'd57320;
ROM1[4242]<=16'd4895; ROM2[4242]<=16'd0; ROM3[4242]<=16'd23804; ROM4[4242]<=16'd57322;
ROM1[4243]<=16'd4858; ROM2[4243]<=16'd0; ROM3[4243]<=16'd23796; ROM4[4243]<=16'd57304;
ROM1[4244]<=16'd4833; ROM2[4244]<=16'd0; ROM3[4244]<=16'd23793; ROM4[4244]<=16'd57293;
ROM1[4245]<=16'd4827; ROM2[4245]<=16'd0; ROM3[4245]<=16'd23801; ROM4[4245]<=16'd57297;
ROM1[4246]<=16'd4816; ROM2[4246]<=16'd0; ROM3[4246]<=16'd23800; ROM4[4246]<=16'd57297;
ROM1[4247]<=16'd4819; ROM2[4247]<=16'd0; ROM3[4247]<=16'd23798; ROM4[4247]<=16'd57298;
ROM1[4248]<=16'd4850; ROM2[4248]<=16'd0; ROM3[4248]<=16'd23792; ROM4[4248]<=16'd57300;
ROM1[4249]<=16'd4887; ROM2[4249]<=16'd0; ROM3[4249]<=16'd23790; ROM4[4249]<=16'd57308;
ROM1[4250]<=16'd4892; ROM2[4250]<=16'd0; ROM3[4250]<=16'd23795; ROM4[4250]<=16'd57313;
ROM1[4251]<=16'd4867; ROM2[4251]<=16'd0; ROM3[4251]<=16'd23792; ROM4[4251]<=16'd57302;
ROM1[4252]<=16'd4853; ROM2[4252]<=16'd0; ROM3[4252]<=16'd23803; ROM4[4252]<=16'd57303;
ROM1[4253]<=16'd4841; ROM2[4253]<=16'd0; ROM3[4253]<=16'd23814; ROM4[4253]<=16'd57304;
ROM1[4254]<=16'd4827; ROM2[4254]<=16'd0; ROM3[4254]<=16'd23824; ROM4[4254]<=16'd57303;
ROM1[4255]<=16'd4837; ROM2[4255]<=16'd0; ROM3[4255]<=16'd23833; ROM4[4255]<=16'd57314;
ROM1[4256]<=16'd4860; ROM2[4256]<=16'd0; ROM3[4256]<=16'd23820; ROM4[4256]<=16'd57311;
ROM1[4257]<=16'd4888; ROM2[4257]<=16'd0; ROM3[4257]<=16'd23802; ROM4[4257]<=16'd57305;
ROM1[4258]<=16'd4900; ROM2[4258]<=16'd0; ROM3[4258]<=16'd23799; ROM4[4258]<=16'd57308;
ROM1[4259]<=16'd4890; ROM2[4259]<=16'd0; ROM3[4259]<=16'd23806; ROM4[4259]<=16'd57311;
ROM1[4260]<=16'd4863; ROM2[4260]<=16'd0; ROM3[4260]<=16'd23807; ROM4[4260]<=16'd57304;
ROM1[4261]<=16'd4846; ROM2[4261]<=16'd0; ROM3[4261]<=16'd23806; ROM4[4261]<=16'd57302;
ROM1[4262]<=16'd4824; ROM2[4262]<=16'd0; ROM3[4262]<=16'd23805; ROM4[4262]<=16'd57297;
ROM1[4263]<=16'd4821; ROM2[4263]<=16'd0; ROM3[4263]<=16'd23810; ROM4[4263]<=16'd57299;
ROM1[4264]<=16'd4859; ROM2[4264]<=16'd0; ROM3[4264]<=16'd23828; ROM4[4264]<=16'd57322;
ROM1[4265]<=16'd4884; ROM2[4265]<=16'd0; ROM3[4265]<=16'd23808; ROM4[4265]<=16'd57314;
ROM1[4266]<=16'd4887; ROM2[4266]<=16'd0; ROM3[4266]<=16'd23780; ROM4[4266]<=16'd57299;
ROM1[4267]<=16'd4876; ROM2[4267]<=16'd0; ROM3[4267]<=16'd23780; ROM4[4267]<=16'd57298;
ROM1[4268]<=16'd4852; ROM2[4268]<=16'd0; ROM3[4268]<=16'd23784; ROM4[4268]<=16'd57293;
ROM1[4269]<=16'd4838; ROM2[4269]<=16'd0; ROM3[4269]<=16'd23796; ROM4[4269]<=16'd57294;
ROM1[4270]<=16'd4829; ROM2[4270]<=16'd0; ROM3[4270]<=16'd23807; ROM4[4270]<=16'd57295;
ROM1[4271]<=16'd4820; ROM2[4271]<=16'd0; ROM3[4271]<=16'd23808; ROM4[4271]<=16'd57296;
ROM1[4272]<=16'd4825; ROM2[4272]<=16'd0; ROM3[4272]<=16'd23803; ROM4[4272]<=16'd57296;
ROM1[4273]<=16'd4855; ROM2[4273]<=16'd0; ROM3[4273]<=16'd23801; ROM4[4273]<=16'd57301;
ROM1[4274]<=16'd4888; ROM2[4274]<=16'd0; ROM3[4274]<=16'd23796; ROM4[4274]<=16'd57306;
ROM1[4275]<=16'd4884; ROM2[4275]<=16'd0; ROM3[4275]<=16'd23796; ROM4[4275]<=16'd57305;
ROM1[4276]<=16'd4863; ROM2[4276]<=16'd0; ROM3[4276]<=16'd23803; ROM4[4276]<=16'd57305;
ROM1[4277]<=16'd4854; ROM2[4277]<=16'd0; ROM3[4277]<=16'd23819; ROM4[4277]<=16'd57316;
ROM1[4278]<=16'd4846; ROM2[4278]<=16'd0; ROM3[4278]<=16'd23827; ROM4[4278]<=16'd57324;
ROM1[4279]<=16'd4847; ROM2[4279]<=16'd0; ROM3[4279]<=16'd23838; ROM4[4279]<=16'd57331;
ROM1[4280]<=16'd4856; ROM2[4280]<=16'd0; ROM3[4280]<=16'd23842; ROM4[4280]<=16'd57337;
ROM1[4281]<=16'd4853; ROM2[4281]<=16'd0; ROM3[4281]<=16'd23808; ROM4[4281]<=16'd57311;
ROM1[4282]<=16'd4873; ROM2[4282]<=16'd0; ROM3[4282]<=16'd23784; ROM4[4282]<=16'd57294;
ROM1[4283]<=16'd4871; ROM2[4283]<=16'd0; ROM3[4283]<=16'd23768; ROM4[4283]<=16'd57284;
ROM1[4284]<=16'd4845; ROM2[4284]<=16'd0; ROM3[4284]<=16'd23757; ROM4[4284]<=16'd57271;
ROM1[4285]<=16'd4838; ROM2[4285]<=16'd0; ROM3[4285]<=16'd23767; ROM4[4285]<=16'd57277;
ROM1[4286]<=16'd4834; ROM2[4286]<=16'd0; ROM3[4286]<=16'd23779; ROM4[4286]<=16'd57281;
ROM1[4287]<=16'd4811; ROM2[4287]<=16'd0; ROM3[4287]<=16'd23775; ROM4[4287]<=16'd57276;
ROM1[4288]<=16'd4798; ROM2[4288]<=16'd0; ROM3[4288]<=16'd23768; ROM4[4288]<=16'd57271;
ROM1[4289]<=16'd4818; ROM2[4289]<=16'd0; ROM3[4289]<=16'd23774; ROM4[4289]<=16'd57281;
ROM1[4290]<=16'd4856; ROM2[4290]<=16'd0; ROM3[4290]<=16'd23774; ROM4[4290]<=16'd57292;
ROM1[4291]<=16'd4887; ROM2[4291]<=16'd0; ROM3[4291]<=16'd23776; ROM4[4291]<=16'd57304;
ROM1[4292]<=16'd4879; ROM2[4292]<=16'd0; ROM3[4292]<=16'd23781; ROM4[4292]<=16'd57306;
ROM1[4293]<=16'd4845; ROM2[4293]<=16'd0; ROM3[4293]<=16'd23774; ROM4[4293]<=16'd57293;
ROM1[4294]<=16'd4820; ROM2[4294]<=16'd0; ROM3[4294]<=16'd23774; ROM4[4294]<=16'd57286;
ROM1[4295]<=16'd4800; ROM2[4295]<=16'd0; ROM3[4295]<=16'd23778; ROM4[4295]<=16'd57280;
ROM1[4296]<=16'd4801; ROM2[4296]<=16'd0; ROM3[4296]<=16'd23789; ROM4[4296]<=16'd57285;
ROM1[4297]<=16'd4820; ROM2[4297]<=16'd0; ROM3[4297]<=16'd23798; ROM4[4297]<=16'd57294;
ROM1[4298]<=16'd4847; ROM2[4298]<=16'd0; ROM3[4298]<=16'd23789; ROM4[4298]<=16'd57297;
ROM1[4299]<=16'd4886; ROM2[4299]<=16'd0; ROM3[4299]<=16'd23787; ROM4[4299]<=16'd57308;
ROM1[4300]<=16'd4888; ROM2[4300]<=16'd0; ROM3[4300]<=16'd23789; ROM4[4300]<=16'd57313;
ROM1[4301]<=16'd4860; ROM2[4301]<=16'd0; ROM3[4301]<=16'd23786; ROM4[4301]<=16'd57307;
ROM1[4302]<=16'd4842; ROM2[4302]<=16'd0; ROM3[4302]<=16'd23794; ROM4[4302]<=16'd57301;
ROM1[4303]<=16'd4826; ROM2[4303]<=16'd0; ROM3[4303]<=16'd23797; ROM4[4303]<=16'd57296;
ROM1[4304]<=16'd4807; ROM2[4304]<=16'd0; ROM3[4304]<=16'd23798; ROM4[4304]<=16'd57288;
ROM1[4305]<=16'd4819; ROM2[4305]<=16'd0; ROM3[4305]<=16'd23807; ROM4[4305]<=16'd57296;
ROM1[4306]<=16'd4847; ROM2[4306]<=16'd0; ROM3[4306]<=16'd23806; ROM4[4306]<=16'd57304;
ROM1[4307]<=16'd4875; ROM2[4307]<=16'd0; ROM3[4307]<=16'd23788; ROM4[4307]<=16'd57297;
ROM1[4308]<=16'd4891; ROM2[4308]<=16'd0; ROM3[4308]<=16'd23787; ROM4[4308]<=16'd57302;
ROM1[4309]<=16'd4874; ROM2[4309]<=16'd0; ROM3[4309]<=16'd23794; ROM4[4309]<=16'd57304;
ROM1[4310]<=16'd4855; ROM2[4310]<=16'd0; ROM3[4310]<=16'd23803; ROM4[4310]<=16'd57304;
ROM1[4311]<=16'd4839; ROM2[4311]<=16'd0; ROM3[4311]<=16'd23807; ROM4[4311]<=16'd57303;
ROM1[4312]<=16'd4805; ROM2[4312]<=16'd0; ROM3[4312]<=16'd23797; ROM4[4312]<=16'd57287;
ROM1[4313]<=16'd4800; ROM2[4313]<=16'd0; ROM3[4313]<=16'd23796; ROM4[4313]<=16'd57285;
ROM1[4314]<=16'd4811; ROM2[4314]<=16'd0; ROM3[4314]<=16'd23788; ROM4[4314]<=16'd57285;
ROM1[4315]<=16'd4831; ROM2[4315]<=16'd0; ROM3[4315]<=16'd23767; ROM4[4315]<=16'd57274;
ROM1[4316]<=16'd4852; ROM2[4316]<=16'd0; ROM3[4316]<=16'd23760; ROM4[4316]<=16'd57271;
ROM1[4317]<=16'd4847; ROM2[4317]<=16'd0; ROM3[4317]<=16'd23763; ROM4[4317]<=16'd57274;
ROM1[4318]<=16'd4828; ROM2[4318]<=16'd0; ROM3[4318]<=16'd23773; ROM4[4318]<=16'd57277;
ROM1[4319]<=16'd4816; ROM2[4319]<=16'd0; ROM3[4319]<=16'd23782; ROM4[4319]<=16'd57276;
ROM1[4320]<=16'd4810; ROM2[4320]<=16'd0; ROM3[4320]<=16'd23794; ROM4[4320]<=16'd57284;
ROM1[4321]<=16'd4803; ROM2[4321]<=16'd0; ROM3[4321]<=16'd23803; ROM4[4321]<=16'd57286;
ROM1[4322]<=16'd4816; ROM2[4322]<=16'd0; ROM3[4322]<=16'd23802; ROM4[4322]<=16'd57287;
ROM1[4323]<=16'd4853; ROM2[4323]<=16'd0; ROM3[4323]<=16'd23798; ROM4[4323]<=16'd57297;
ROM1[4324]<=16'd4886; ROM2[4324]<=16'd0; ROM3[4324]<=16'd23792; ROM4[4324]<=16'd57305;
ROM1[4325]<=16'd4889; ROM2[4325]<=16'd0; ROM3[4325]<=16'd23790; ROM4[4325]<=16'd57306;
ROM1[4326]<=16'd4868; ROM2[4326]<=16'd0; ROM3[4326]<=16'd23790; ROM4[4326]<=16'd57301;
ROM1[4327]<=16'd4845; ROM2[4327]<=16'd0; ROM3[4327]<=16'd23799; ROM4[4327]<=16'd57300;
ROM1[4328]<=16'd4832; ROM2[4328]<=16'd0; ROM3[4328]<=16'd23805; ROM4[4328]<=16'd57301;
ROM1[4329]<=16'd4818; ROM2[4329]<=16'd0; ROM3[4329]<=16'd23806; ROM4[4329]<=16'd57297;
ROM1[4330]<=16'd4825; ROM2[4330]<=16'd0; ROM3[4330]<=16'd23810; ROM4[4330]<=16'd57301;
ROM1[4331]<=16'd4866; ROM2[4331]<=16'd0; ROM3[4331]<=16'd23824; ROM4[4331]<=16'd57320;
ROM1[4332]<=16'd4905; ROM2[4332]<=16'd0; ROM3[4332]<=16'd23819; ROM4[4332]<=16'd57324;
ROM1[4333]<=16'd4892; ROM2[4333]<=16'd0; ROM3[4333]<=16'd23797; ROM4[4333]<=16'd57306;
ROM1[4334]<=16'd4867; ROM2[4334]<=16'd0; ROM3[4334]<=16'd23794; ROM4[4334]<=16'd57298;
ROM1[4335]<=16'd4833; ROM2[4335]<=16'd0; ROM3[4335]<=16'd23780; ROM4[4335]<=16'd57281;
ROM1[4336]<=16'd4821; ROM2[4336]<=16'd0; ROM3[4336]<=16'd23785; ROM4[4336]<=16'd57282;
ROM1[4337]<=16'd4820; ROM2[4337]<=16'd0; ROM3[4337]<=16'd23807; ROM4[4337]<=16'd57297;
ROM1[4338]<=16'd4807; ROM2[4338]<=16'd0; ROM3[4338]<=16'd23801; ROM4[4338]<=16'd57289;
ROM1[4339]<=16'd4817; ROM2[4339]<=16'd0; ROM3[4339]<=16'd23789; ROM4[4339]<=16'd57281;
ROM1[4340]<=16'd4849; ROM2[4340]<=16'd0; ROM3[4340]<=16'd23778; ROM4[4340]<=16'd57284;
ROM1[4341]<=16'd4886; ROM2[4341]<=16'd0; ROM3[4341]<=16'd23783; ROM4[4341]<=16'd57298;
ROM1[4342]<=16'd4889; ROM2[4342]<=16'd0; ROM3[4342]<=16'd23792; ROM4[4342]<=16'd57305;
ROM1[4343]<=16'd4867; ROM2[4343]<=16'd0; ROM3[4343]<=16'd23791; ROM4[4343]<=16'd57299;
ROM1[4344]<=16'd4843; ROM2[4344]<=16'd0; ROM3[4344]<=16'd23789; ROM4[4344]<=16'd57290;
ROM1[4345]<=16'd4825; ROM2[4345]<=16'd0; ROM3[4345]<=16'd23786; ROM4[4345]<=16'd57283;
ROM1[4346]<=16'd4811; ROM2[4346]<=16'd0; ROM3[4346]<=16'd23788; ROM4[4346]<=16'd57278;
ROM1[4347]<=16'd4814; ROM2[4347]<=16'd0; ROM3[4347]<=16'd23788; ROM4[4347]<=16'd57274;
ROM1[4348]<=16'd4845; ROM2[4348]<=16'd0; ROM3[4348]<=16'd23783; ROM4[4348]<=16'd57275;
ROM1[4349]<=16'd4872; ROM2[4349]<=16'd0; ROM3[4349]<=16'd23768; ROM4[4349]<=16'd57274;
ROM1[4350]<=16'd4871; ROM2[4350]<=16'd0; ROM3[4350]<=16'd23765; ROM4[4350]<=16'd57274;
ROM1[4351]<=16'd4857; ROM2[4351]<=16'd0; ROM3[4351]<=16'd23779; ROM4[4351]<=16'd57278;
ROM1[4352]<=16'd4839; ROM2[4352]<=16'd0; ROM3[4352]<=16'd23788; ROM4[4352]<=16'd57280;
ROM1[4353]<=16'd4821; ROM2[4353]<=16'd0; ROM3[4353]<=16'd23792; ROM4[4353]<=16'd57278;
ROM1[4354]<=16'd4812; ROM2[4354]<=16'd0; ROM3[4354]<=16'd23804; ROM4[4354]<=16'd57283;
ROM1[4355]<=16'd4819; ROM2[4355]<=16'd0; ROM3[4355]<=16'd23806; ROM4[4355]<=16'd57286;
ROM1[4356]<=16'd4836; ROM2[4356]<=16'd0; ROM3[4356]<=16'd23793; ROM4[4356]<=16'd57282;
ROM1[4357]<=16'd4865; ROM2[4357]<=16'd0; ROM3[4357]<=16'd23777; ROM4[4357]<=16'd57278;
ROM1[4358]<=16'd4872; ROM2[4358]<=16'd0; ROM3[4358]<=16'd23769; ROM4[4358]<=16'd57271;
ROM1[4359]<=16'd4860; ROM2[4359]<=16'd0; ROM3[4359]<=16'd23774; ROM4[4359]<=16'd57272;
ROM1[4360]<=16'd4851; ROM2[4360]<=16'd0; ROM3[4360]<=16'd23787; ROM4[4360]<=16'd57280;
ROM1[4361]<=16'd4859; ROM2[4361]<=16'd0; ROM3[4361]<=16'd23811; ROM4[4361]<=16'd57301;
ROM1[4362]<=16'd4849; ROM2[4362]<=16'd0; ROM3[4362]<=16'd23819; ROM4[4362]<=16'd57306;
ROM1[4363]<=16'd4828; ROM2[4363]<=16'd0; ROM3[4363]<=16'd23805; ROM4[4363]<=16'd57288;
ROM1[4364]<=16'd4839; ROM2[4364]<=16'd0; ROM3[4364]<=16'd23800; ROM4[4364]<=16'd57289;
ROM1[4365]<=16'd4866; ROM2[4365]<=16'd0; ROM3[4365]<=16'd23785; ROM4[4365]<=16'd57288;
ROM1[4366]<=16'd4878; ROM2[4366]<=16'd0; ROM3[4366]<=16'd23773; ROM4[4366]<=16'd57284;
ROM1[4367]<=16'd4880; ROM2[4367]<=16'd0; ROM3[4367]<=16'd23786; ROM4[4367]<=16'd57293;
ROM1[4368]<=16'd4872; ROM2[4368]<=16'd0; ROM3[4368]<=16'd23807; ROM4[4368]<=16'd57303;
ROM1[4369]<=16'd4855; ROM2[4369]<=16'd0; ROM3[4369]<=16'd23815; ROM4[4369]<=16'd57301;
ROM1[4370]<=16'd4841; ROM2[4370]<=16'd0; ROM3[4370]<=16'd23819; ROM4[4370]<=16'd57301;
ROM1[4371]<=16'd4834; ROM2[4371]<=16'd0; ROM3[4371]<=16'd23829; ROM4[4371]<=16'd57309;
ROM1[4372]<=16'd4836; ROM2[4372]<=16'd0; ROM3[4372]<=16'd23823; ROM4[4372]<=16'd57304;
ROM1[4373]<=16'd4862; ROM2[4373]<=16'd0; ROM3[4373]<=16'd23808; ROM4[4373]<=16'd57298;
ROM1[4374]<=16'd4892; ROM2[4374]<=16'd0; ROM3[4374]<=16'd23799; ROM4[4374]<=16'd57300;
ROM1[4375]<=16'd4883; ROM2[4375]<=16'd0; ROM3[4375]<=16'd23790; ROM4[4375]<=16'd57294;
ROM1[4376]<=16'd4857; ROM2[4376]<=16'd0; ROM3[4376]<=16'd23783; ROM4[4376]<=16'd57284;
ROM1[4377]<=16'd4840; ROM2[4377]<=16'd0; ROM3[4377]<=16'd23791; ROM4[4377]<=16'd57285;
ROM1[4378]<=16'd4830; ROM2[4378]<=16'd0; ROM3[4378]<=16'd23798; ROM4[4378]<=16'd57290;
ROM1[4379]<=16'd4822; ROM2[4379]<=16'd0; ROM3[4379]<=16'd23804; ROM4[4379]<=16'd57291;
ROM1[4380]<=16'd4826; ROM2[4380]<=16'd0; ROM3[4380]<=16'd23804; ROM4[4380]<=16'd57293;
ROM1[4381]<=16'd4846; ROM2[4381]<=16'd0; ROM3[4381]<=16'd23797; ROM4[4381]<=16'd57294;
ROM1[4382]<=16'd4878; ROM2[4382]<=16'd0; ROM3[4382]<=16'd23785; ROM4[4382]<=16'd57295;
ROM1[4383]<=16'd4900; ROM2[4383]<=16'd0; ROM3[4383]<=16'd23782; ROM4[4383]<=16'd57305;
ROM1[4384]<=16'd4899; ROM2[4384]<=16'd0; ROM3[4384]<=16'd23792; ROM4[4384]<=16'd57312;
ROM1[4385]<=16'd4883; ROM2[4385]<=16'd0; ROM3[4385]<=16'd23802; ROM4[4385]<=16'd57312;
ROM1[4386]<=16'd4862; ROM2[4386]<=16'd0; ROM3[4386]<=16'd23796; ROM4[4386]<=16'd57304;
ROM1[4387]<=16'd4824; ROM2[4387]<=16'd0; ROM3[4387]<=16'd23780; ROM4[4387]<=16'd57281;
ROM1[4388]<=16'd4812; ROM2[4388]<=16'd0; ROM3[4388]<=16'd23775; ROM4[4388]<=16'd57276;
ROM1[4389]<=16'd4831; ROM2[4389]<=16'd0; ROM3[4389]<=16'd23776; ROM4[4389]<=16'd57284;
ROM1[4390]<=16'd4871; ROM2[4390]<=16'd0; ROM3[4390]<=16'd23773; ROM4[4390]<=16'd57287;
ROM1[4391]<=16'd4893; ROM2[4391]<=16'd0; ROM3[4391]<=16'd23772; ROM4[4391]<=16'd57296;
ROM1[4392]<=16'd4875; ROM2[4392]<=16'd0; ROM3[4392]<=16'd23765; ROM4[4392]<=16'd57289;
ROM1[4393]<=16'd4847; ROM2[4393]<=16'd0; ROM3[4393]<=16'd23758; ROM4[4393]<=16'd57275;
ROM1[4394]<=16'd4832; ROM2[4394]<=16'd0; ROM3[4394]<=16'd23767; ROM4[4394]<=16'd57278;
ROM1[4395]<=16'd4823; ROM2[4395]<=16'd0; ROM3[4395]<=16'd23776; ROM4[4395]<=16'd57279;
ROM1[4396]<=16'd4815; ROM2[4396]<=16'd0; ROM3[4396]<=16'd23782; ROM4[4396]<=16'd57280;
ROM1[4397]<=16'd4828; ROM2[4397]<=16'd0; ROM3[4397]<=16'd23786; ROM4[4397]<=16'd57286;
ROM1[4398]<=16'd4859; ROM2[4398]<=16'd0; ROM3[4398]<=16'd23778; ROM4[4398]<=16'd57288;
ROM1[4399]<=16'd4892; ROM2[4399]<=16'd0; ROM3[4399]<=16'd23775; ROM4[4399]<=16'd57294;
ROM1[4400]<=16'd4895; ROM2[4400]<=16'd0; ROM3[4400]<=16'd23782; ROM4[4400]<=16'd57300;
ROM1[4401]<=16'd4875; ROM2[4401]<=16'd0; ROM3[4401]<=16'd23792; ROM4[4401]<=16'd57302;
ROM1[4402]<=16'd4852; ROM2[4402]<=16'd0; ROM3[4402]<=16'd23800; ROM4[4402]<=16'd57298;
ROM1[4403]<=16'd4847; ROM2[4403]<=16'd0; ROM3[4403]<=16'd23813; ROM4[4403]<=16'd57304;
ROM1[4404]<=16'd4843; ROM2[4404]<=16'd0; ROM3[4404]<=16'd23819; ROM4[4404]<=16'd57306;
ROM1[4405]<=16'd4827; ROM2[4405]<=16'd0; ROM3[4405]<=16'd23800; ROM4[4405]<=16'd57286;
ROM1[4406]<=16'd4829; ROM2[4406]<=16'd0; ROM3[4406]<=16'd23772; ROM4[4406]<=16'd57270;
ROM1[4407]<=16'd4859; ROM2[4407]<=16'd0; ROM3[4407]<=16'd23754; ROM4[4407]<=16'd57269;
ROM1[4408]<=16'd4866; ROM2[4408]<=16'd0; ROM3[4408]<=16'd23751; ROM4[4408]<=16'd57269;
ROM1[4409]<=16'd4853; ROM2[4409]<=16'd0; ROM3[4409]<=16'd23756; ROM4[4409]<=16'd57271;
ROM1[4410]<=16'd4847; ROM2[4410]<=16'd0; ROM3[4410]<=16'd23772; ROM4[4410]<=16'd57281;
ROM1[4411]<=16'd4834; ROM2[4411]<=16'd0; ROM3[4411]<=16'd23786; ROM4[4411]<=16'd57289;
ROM1[4412]<=16'd4810; ROM2[4412]<=16'd0; ROM3[4412]<=16'd23784; ROM4[4412]<=16'd57284;
ROM1[4413]<=16'd4809; ROM2[4413]<=16'd0; ROM3[4413]<=16'd23785; ROM4[4413]<=16'd57282;
ROM1[4414]<=16'd4823; ROM2[4414]<=16'd0; ROM3[4414]<=16'd23779; ROM4[4414]<=16'd57279;
ROM1[4415]<=16'd4857; ROM2[4415]<=16'd0; ROM3[4415]<=16'd23773; ROM4[4415]<=16'd57282;
ROM1[4416]<=16'd4894; ROM2[4416]<=16'd0; ROM3[4416]<=16'd23785; ROM4[4416]<=16'd57297;
ROM1[4417]<=16'd4896; ROM2[4417]<=16'd0; ROM3[4417]<=16'd23799; ROM4[4417]<=16'd57313;
ROM1[4418]<=16'd4874; ROM2[4418]<=16'd0; ROM3[4418]<=16'd23803; ROM4[4418]<=16'd57310;
ROM1[4419]<=16'd4857; ROM2[4419]<=16'd0; ROM3[4419]<=16'd23806; ROM4[4419]<=16'd57305;
ROM1[4420]<=16'd4831; ROM2[4420]<=16'd0; ROM3[4420]<=16'd23800; ROM4[4420]<=16'd57295;
ROM1[4421]<=16'd4811; ROM2[4421]<=16'd0; ROM3[4421]<=16'd23796; ROM4[4421]<=16'd57283;
ROM1[4422]<=16'd4827; ROM2[4422]<=16'd0; ROM3[4422]<=16'd23803; ROM4[4422]<=16'd57293;
ROM1[4423]<=16'd4848; ROM2[4423]<=16'd0; ROM3[4423]<=16'd23789; ROM4[4423]<=16'd57286;
ROM1[4424]<=16'd4871; ROM2[4424]<=16'd0; ROM3[4424]<=16'd23775; ROM4[4424]<=16'd57282;
ROM1[4425]<=16'd4872; ROM2[4425]<=16'd0; ROM3[4425]<=16'd23773; ROM4[4425]<=16'd57285;
ROM1[4426]<=16'd4854; ROM2[4426]<=16'd0; ROM3[4426]<=16'd23775; ROM4[4426]<=16'd57282;
ROM1[4427]<=16'd4831; ROM2[4427]<=16'd0; ROM3[4427]<=16'd23779; ROM4[4427]<=16'd57281;
ROM1[4428]<=16'd4817; ROM2[4428]<=16'd0; ROM3[4428]<=16'd23784; ROM4[4428]<=16'd57278;
ROM1[4429]<=16'd4805; ROM2[4429]<=16'd0; ROM3[4429]<=16'd23787; ROM4[4429]<=16'd57273;
ROM1[4430]<=16'd4800; ROM2[4430]<=16'd0; ROM3[4430]<=16'd23780; ROM4[4430]<=16'd57267;
ROM1[4431]<=16'd4827; ROM2[4431]<=16'd0; ROM3[4431]<=16'd23770; ROM4[4431]<=16'd57267;
ROM1[4432]<=16'd4868; ROM2[4432]<=16'd0; ROM3[4432]<=16'd23763; ROM4[4432]<=16'd57272;
ROM1[4433]<=16'd4873; ROM2[4433]<=16'd0; ROM3[4433]<=16'd23759; ROM4[4433]<=16'd57271;
ROM1[4434]<=16'd4865; ROM2[4434]<=16'd0; ROM3[4434]<=16'd23765; ROM4[4434]<=16'd57271;
ROM1[4435]<=16'd4856; ROM2[4435]<=16'd0; ROM3[4435]<=16'd23779; ROM4[4435]<=16'd57275;
ROM1[4436]<=16'd4837; ROM2[4436]<=16'd0; ROM3[4436]<=16'd23778; ROM4[4436]<=16'd57271;
ROM1[4437]<=16'd4822; ROM2[4437]<=16'd0; ROM3[4437]<=16'd23784; ROM4[4437]<=16'd57275;
ROM1[4438]<=16'd4842; ROM2[4438]<=16'd0; ROM3[4438]<=16'd23807; ROM4[4438]<=16'd57298;
ROM1[4439]<=16'd4842; ROM2[4439]<=16'd0; ROM3[4439]<=16'd23790; ROM4[4439]<=16'd57288;
ROM1[4440]<=16'd4840; ROM2[4440]<=16'd0; ROM3[4440]<=16'd23749; ROM4[4440]<=16'd57256;
ROM1[4441]<=16'd4864; ROM2[4441]<=16'd0; ROM3[4441]<=16'd23745; ROM4[4441]<=16'd57264;
ROM1[4442]<=16'd4858; ROM2[4442]<=16'd0; ROM3[4442]<=16'd23753; ROM4[4442]<=16'd57269;
ROM1[4443]<=16'd4853; ROM2[4443]<=16'd0; ROM3[4443]<=16'd23767; ROM4[4443]<=16'd57277;
ROM1[4444]<=16'd4855; ROM2[4444]<=16'd0; ROM3[4444]<=16'd23787; ROM4[4444]<=16'd57292;
ROM1[4445]<=16'd4828; ROM2[4445]<=16'd0; ROM3[4445]<=16'd23779; ROM4[4445]<=16'd57278;
ROM1[4446]<=16'd4808; ROM2[4446]<=16'd0; ROM3[4446]<=16'd23773; ROM4[4446]<=16'd57267;
ROM1[4447]<=16'd4811; ROM2[4447]<=16'd0; ROM3[4447]<=16'd23766; ROM4[4447]<=16'd57264;
ROM1[4448]<=16'd4841; ROM2[4448]<=16'd0; ROM3[4448]<=16'd23761; ROM4[4448]<=16'd57267;
ROM1[4449]<=16'd4879; ROM2[4449]<=16'd0; ROM3[4449]<=16'd23760; ROM4[4449]<=16'd57275;
ROM1[4450]<=16'd4881; ROM2[4450]<=16'd0; ROM3[4450]<=16'd23763; ROM4[4450]<=16'd57277;
ROM1[4451]<=16'd4872; ROM2[4451]<=16'd0; ROM3[4451]<=16'd23778; ROM4[4451]<=16'd57287;
ROM1[4452]<=16'd4857; ROM2[4452]<=16'd0; ROM3[4452]<=16'd23787; ROM4[4452]<=16'd57290;
ROM1[4453]<=16'd4829; ROM2[4453]<=16'd0; ROM3[4453]<=16'd23778; ROM4[4453]<=16'd57276;
ROM1[4454]<=16'd4804; ROM2[4454]<=16'd0; ROM3[4454]<=16'd23768; ROM4[4454]<=16'd57261;
ROM1[4455]<=16'd4803; ROM2[4455]<=16'd0; ROM3[4455]<=16'd23765; ROM4[4455]<=16'd57255;
ROM1[4456]<=16'd4819; ROM2[4456]<=16'd0; ROM3[4456]<=16'd23755; ROM4[4456]<=16'd57250;
ROM1[4457]<=16'd4864; ROM2[4457]<=16'd0; ROM3[4457]<=16'd23755; ROM4[4457]<=16'd57261;
ROM1[4458]<=16'd4877; ROM2[4458]<=16'd0; ROM3[4458]<=16'd23754; ROM4[4458]<=16'd57266;
ROM1[4459]<=16'd4858; ROM2[4459]<=16'd0; ROM3[4459]<=16'd23749; ROM4[4459]<=16'd57263;
ROM1[4460]<=16'd4849; ROM2[4460]<=16'd0; ROM3[4460]<=16'd23761; ROM4[4460]<=16'd57270;
ROM1[4461]<=16'd4839; ROM2[4461]<=16'd0; ROM3[4461]<=16'd23769; ROM4[4461]<=16'd57268;
ROM1[4462]<=16'd4836; ROM2[4462]<=16'd0; ROM3[4462]<=16'd23786; ROM4[4462]<=16'd57282;
ROM1[4463]<=16'd4841; ROM2[4463]<=16'd0; ROM3[4463]<=16'd23800; ROM4[4463]<=16'd57291;
ROM1[4464]<=16'd4855; ROM2[4464]<=16'd0; ROM3[4464]<=16'd23797; ROM4[4464]<=16'd57287;
ROM1[4465]<=16'd4882; ROM2[4465]<=16'd0; ROM3[4465]<=16'd23783; ROM4[4465]<=16'd57287;
ROM1[4466]<=16'd4892; ROM2[4466]<=16'd0; ROM3[4466]<=16'd23766; ROM4[4466]<=16'd57278;
ROM1[4467]<=16'd4883; ROM2[4467]<=16'd0; ROM3[4467]<=16'd23767; ROM4[4467]<=16'd57276;
ROM1[4468]<=16'd4862; ROM2[4468]<=16'd0; ROM3[4468]<=16'd23776; ROM4[4468]<=16'd57276;
ROM1[4469]<=16'd4851; ROM2[4469]<=16'd0; ROM3[4469]<=16'd23785; ROM4[4469]<=16'd57280;
ROM1[4470]<=16'd4833; ROM2[4470]<=16'd0; ROM3[4470]<=16'd23788; ROM4[4470]<=16'd57281;
ROM1[4471]<=16'd4813; ROM2[4471]<=16'd0; ROM3[4471]<=16'd23784; ROM4[4471]<=16'd57271;
ROM1[4472]<=16'd4827; ROM2[4472]<=16'd0; ROM3[4472]<=16'd23785; ROM4[4472]<=16'd57276;
ROM1[4473]<=16'd4864; ROM2[4473]<=16'd0; ROM3[4473]<=16'd23786; ROM4[4473]<=16'd57289;
ROM1[4474]<=16'd4886; ROM2[4474]<=16'd0; ROM3[4474]<=16'd23772; ROM4[4474]<=16'd57284;
ROM1[4475]<=16'd4879; ROM2[4475]<=16'd0; ROM3[4475]<=16'd23772; ROM4[4475]<=16'd57280;
ROM1[4476]<=16'd4867; ROM2[4476]<=16'd0; ROM3[4476]<=16'd23789; ROM4[4476]<=16'd57288;
ROM1[4477]<=16'd4853; ROM2[4477]<=16'd0; ROM3[4477]<=16'd23798; ROM4[4477]<=16'd57288;
ROM1[4478]<=16'd4836; ROM2[4478]<=16'd0; ROM3[4478]<=16'd23803; ROM4[4478]<=16'd57285;
ROM1[4479]<=16'd4823; ROM2[4479]<=16'd0; ROM3[4479]<=16'd23810; ROM4[4479]<=16'd57284;
ROM1[4480]<=16'd4829; ROM2[4480]<=16'd0; ROM3[4480]<=16'd23813; ROM4[4480]<=16'd57287;
ROM1[4481]<=16'd4845; ROM2[4481]<=16'd0; ROM3[4481]<=16'd23803; ROM4[4481]<=16'd57284;
ROM1[4482]<=16'd4874; ROM2[4482]<=16'd0; ROM3[4482]<=16'd23790; ROM4[4482]<=16'd57281;
ROM1[4483]<=16'd4886; ROM2[4483]<=16'd0; ROM3[4483]<=16'd23788; ROM4[4483]<=16'd57282;
ROM1[4484]<=16'd4874; ROM2[4484]<=16'd0; ROM3[4484]<=16'd23790; ROM4[4484]<=16'd57280;
ROM1[4485]<=16'd4852; ROM2[4485]<=16'd0; ROM3[4485]<=16'd23793; ROM4[4485]<=16'd57273;
ROM1[4486]<=16'd4839; ROM2[4486]<=16'd0; ROM3[4486]<=16'd23798; ROM4[4486]<=16'd57274;
ROM1[4487]<=16'd4826; ROM2[4487]<=16'd0; ROM3[4487]<=16'd23806; ROM4[4487]<=16'd57281;
ROM1[4488]<=16'd4818; ROM2[4488]<=16'd0; ROM3[4488]<=16'd23803; ROM4[4488]<=16'd57280;
ROM1[4489]<=16'd4845; ROM2[4489]<=16'd0; ROM3[4489]<=16'd23808; ROM4[4489]<=16'd57291;
ROM1[4490]<=16'd4890; ROM2[4490]<=16'd0; ROM3[4490]<=16'd23812; ROM4[4490]<=16'd57302;
ROM1[4491]<=16'd4884; ROM2[4491]<=16'd0; ROM3[4491]<=16'd23778; ROM4[4491]<=16'd57275;
ROM1[4492]<=16'd4862; ROM2[4492]<=16'd0; ROM3[4492]<=16'd23765; ROM4[4492]<=16'd57262;
ROM1[4493]<=16'd4844; ROM2[4493]<=16'd0; ROM3[4493]<=16'd23773; ROM4[4493]<=16'd57263;
ROM1[4494]<=16'd4826; ROM2[4494]<=16'd0; ROM3[4494]<=16'd23783; ROM4[4494]<=16'd57266;
ROM1[4495]<=16'd4831; ROM2[4495]<=16'd0; ROM3[4495]<=16'd23809; ROM4[4495]<=16'd57290;
ROM1[4496]<=16'd4838; ROM2[4496]<=16'd0; ROM3[4496]<=16'd23824; ROM4[4496]<=16'd57302;
ROM1[4497]<=16'd4835; ROM2[4497]<=16'd0; ROM3[4497]<=16'd23809; ROM4[4497]<=16'd57292;
ROM1[4498]<=16'd4857; ROM2[4498]<=16'd0; ROM3[4498]<=16'd23789; ROM4[4498]<=16'd57288;
ROM1[4499]<=16'd4901; ROM2[4499]<=16'd0; ROM3[4499]<=16'd23790; ROM4[4499]<=16'd57303;
ROM1[4500]<=16'd4897; ROM2[4500]<=16'd0; ROM3[4500]<=16'd23788; ROM4[4500]<=16'd57302;
ROM1[4501]<=16'd4882; ROM2[4501]<=16'd0; ROM3[4501]<=16'd23800; ROM4[4501]<=16'd57309;
ROM1[4502]<=16'd4872; ROM2[4502]<=16'd0; ROM3[4502]<=16'd23821; ROM4[4502]<=16'd57319;
ROM1[4503]<=16'd4833; ROM2[4503]<=16'd0; ROM3[4503]<=16'd23805; ROM4[4503]<=16'd57298;
ROM1[4504]<=16'd4810; ROM2[4504]<=16'd0; ROM3[4504]<=16'd23802; ROM4[4504]<=16'd57293;
ROM1[4505]<=16'd4814; ROM2[4505]<=16'd0; ROM3[4505]<=16'd23801; ROM4[4505]<=16'd57290;
ROM1[4506]<=16'd4830; ROM2[4506]<=16'd0; ROM3[4506]<=16'd23781; ROM4[4506]<=16'd57275;
ROM1[4507]<=16'd4877; ROM2[4507]<=16'd0; ROM3[4507]<=16'd23777; ROM4[4507]<=16'd57281;
ROM1[4508]<=16'd4895; ROM2[4508]<=16'd0; ROM3[4508]<=16'd23786; ROM4[4508]<=16'd57292;
ROM1[4509]<=16'd4883; ROM2[4509]<=16'd0; ROM3[4509]<=16'd23794; ROM4[4509]<=16'd57296;
ROM1[4510]<=16'd4863; ROM2[4510]<=16'd0; ROM3[4510]<=16'd23799; ROM4[4510]<=16'd57295;
ROM1[4511]<=16'd4852; ROM2[4511]<=16'd0; ROM3[4511]<=16'd23810; ROM4[4511]<=16'd57299;
ROM1[4512]<=16'd4836; ROM2[4512]<=16'd0; ROM3[4512]<=16'd23813; ROM4[4512]<=16'd57298;
ROM1[4513]<=16'd4825; ROM2[4513]<=16'd0; ROM3[4513]<=16'd23806; ROM4[4513]<=16'd57288;
ROM1[4514]<=16'd4839; ROM2[4514]<=16'd0; ROM3[4514]<=16'd23796; ROM4[4514]<=16'd57282;
ROM1[4515]<=16'd4870; ROM2[4515]<=16'd0; ROM3[4515]<=16'd23782; ROM4[4515]<=16'd57285;
ROM1[4516]<=16'd4890; ROM2[4516]<=16'd0; ROM3[4516]<=16'd23775; ROM4[4516]<=16'd57286;
ROM1[4517]<=16'd4879; ROM2[4517]<=16'd0; ROM3[4517]<=16'd23780; ROM4[4517]<=16'd57286;
ROM1[4518]<=16'd4867; ROM2[4518]<=16'd0; ROM3[4518]<=16'd23791; ROM4[4518]<=16'd57293;
ROM1[4519]<=16'd4860; ROM2[4519]<=16'd0; ROM3[4519]<=16'd23805; ROM4[4519]<=16'd57300;
ROM1[4520]<=16'd4855; ROM2[4520]<=16'd0; ROM3[4520]<=16'd23816; ROM4[4520]<=16'd57305;
ROM1[4521]<=16'd4843; ROM2[4521]<=16'd0; ROM3[4521]<=16'd23814; ROM4[4521]<=16'd57303;
ROM1[4522]<=16'd4846; ROM2[4522]<=16'd0; ROM3[4522]<=16'd23805; ROM4[4522]<=16'd57298;
ROM1[4523]<=16'd4879; ROM2[4523]<=16'd0; ROM3[4523]<=16'd23802; ROM4[4523]<=16'd57300;
ROM1[4524]<=16'd4910; ROM2[4524]<=16'd0; ROM3[4524]<=16'd23800; ROM4[4524]<=16'd57307;
ROM1[4525]<=16'd4902; ROM2[4525]<=16'd0; ROM3[4525]<=16'd23798; ROM4[4525]<=16'd57303;
ROM1[4526]<=16'd4887; ROM2[4526]<=16'd0; ROM3[4526]<=16'd23810; ROM4[4526]<=16'd57309;
ROM1[4527]<=16'd4865; ROM2[4527]<=16'd0; ROM3[4527]<=16'd23815; ROM4[4527]<=16'd57305;
ROM1[4528]<=16'd4834; ROM2[4528]<=16'd0; ROM3[4528]<=16'd23808; ROM4[4528]<=16'd57291;
ROM1[4529]<=16'd4823; ROM2[4529]<=16'd0; ROM3[4529]<=16'd23815; ROM4[4529]<=16'd57296;
ROM1[4530]<=16'd4826; ROM2[4530]<=16'd0; ROM3[4530]<=16'd23814; ROM4[4530]<=16'd57294;
ROM1[4531]<=16'd4841; ROM2[4531]<=16'd0; ROM3[4531]<=16'd23794; ROM4[4531]<=16'd57285;
ROM1[4532]<=16'd4871; ROM2[4532]<=16'd0; ROM3[4532]<=16'd23778; ROM4[4532]<=16'd57280;
ROM1[4533]<=16'd4883; ROM2[4533]<=16'd0; ROM3[4533]<=16'd23779; ROM4[4533]<=16'd57285;
ROM1[4534]<=16'd4868; ROM2[4534]<=16'd0; ROM3[4534]<=16'd23782; ROM4[4534]<=16'd57287;
ROM1[4535]<=16'd4853; ROM2[4535]<=16'd0; ROM3[4535]<=16'd23796; ROM4[4535]<=16'd57295;
ROM1[4536]<=16'd4856; ROM2[4536]<=16'd0; ROM3[4536]<=16'd23821; ROM4[4536]<=16'd57316;
ROM1[4537]<=16'd4842; ROM2[4537]<=16'd0; ROM3[4537]<=16'd23825; ROM4[4537]<=16'd57312;
ROM1[4538]<=16'd4829; ROM2[4538]<=16'd0; ROM3[4538]<=16'd23814; ROM4[4538]<=16'd57296;
ROM1[4539]<=16'd4837; ROM2[4539]<=16'd0; ROM3[4539]<=16'd23801; ROM4[4539]<=16'd57286;
ROM1[4540]<=16'd4844; ROM2[4540]<=16'd0; ROM3[4540]<=16'd23767; ROM4[4540]<=16'd57264;
ROM1[4541]<=16'd4857; ROM2[4541]<=16'd0; ROM3[4541]<=16'd23753; ROM4[4541]<=16'd57257;
ROM1[4542]<=16'd4854; ROM2[4542]<=16'd0; ROM3[4542]<=16'd23771; ROM4[4542]<=16'd57269;
ROM1[4543]<=16'd4839; ROM2[4543]<=16'd0; ROM3[4543]<=16'd23784; ROM4[4543]<=16'd57275;
ROM1[4544]<=16'd4825; ROM2[4544]<=16'd0; ROM3[4544]<=16'd23792; ROM4[4544]<=16'd57273;
ROM1[4545]<=16'd4806; ROM2[4545]<=16'd0; ROM3[4545]<=16'd23794; ROM4[4545]<=16'd57271;
ROM1[4546]<=16'd4798; ROM2[4546]<=16'd0; ROM3[4546]<=16'd23797; ROM4[4546]<=16'd57276;
ROM1[4547]<=16'd4805; ROM2[4547]<=16'd0; ROM3[4547]<=16'd23790; ROM4[4547]<=16'd57271;
ROM1[4548]<=16'd4830; ROM2[4548]<=16'd0; ROM3[4548]<=16'd23773; ROM4[4548]<=16'd57268;
ROM1[4549]<=16'd4858; ROM2[4549]<=16'd0; ROM3[4549]<=16'd23759; ROM4[4549]<=16'd57271;
ROM1[4550]<=16'd4853; ROM2[4550]<=16'd0; ROM3[4550]<=16'd23750; ROM4[4550]<=16'd57265;
ROM1[4551]<=16'd4828; ROM2[4551]<=16'd0; ROM3[4551]<=16'd23745; ROM4[4551]<=16'd57255;
ROM1[4552]<=16'd4825; ROM2[4552]<=16'd0; ROM3[4552]<=16'd23760; ROM4[4552]<=16'd57265;
ROM1[4553]<=16'd4835; ROM2[4553]<=16'd0; ROM3[4553]<=16'd23785; ROM4[4553]<=16'd57282;
ROM1[4554]<=16'd4811; ROM2[4554]<=16'd0; ROM3[4554]<=16'd23778; ROM4[4554]<=16'd57272;
ROM1[4555]<=16'd4797; ROM2[4555]<=16'd0; ROM3[4555]<=16'd23760; ROM4[4555]<=16'd57258;
ROM1[4556]<=16'd4816; ROM2[4556]<=16'd0; ROM3[4556]<=16'd23752; ROM4[4556]<=16'd57250;
ROM1[4557]<=16'd4842; ROM2[4557]<=16'd0; ROM3[4557]<=16'd23737; ROM4[4557]<=16'd57245;
ROM1[4558]<=16'd4854; ROM2[4558]<=16'd0; ROM3[4558]<=16'd23738; ROM4[4558]<=16'd57247;
ROM1[4559]<=16'd4853; ROM2[4559]<=16'd0; ROM3[4559]<=16'd23758; ROM4[4559]<=16'd57261;
ROM1[4560]<=16'd4831; ROM2[4560]<=16'd0; ROM3[4560]<=16'd23763; ROM4[4560]<=16'd57262;
ROM1[4561]<=16'd4814; ROM2[4561]<=16'd0; ROM3[4561]<=16'd23764; ROM4[4561]<=16'd57258;
ROM1[4562]<=16'd4810; ROM2[4562]<=16'd0; ROM3[4562]<=16'd23778; ROM4[4562]<=16'd57268;
ROM1[4563]<=16'd4813; ROM2[4563]<=16'd0; ROM3[4563]<=16'd23789; ROM4[4563]<=16'd57276;
ROM1[4564]<=16'd4820; ROM2[4564]<=16'd0; ROM3[4564]<=16'd23779; ROM4[4564]<=16'd57269;
ROM1[4565]<=16'd4847; ROM2[4565]<=16'd0; ROM3[4565]<=16'd23766; ROM4[4565]<=16'd57266;
ROM1[4566]<=16'd4875; ROM2[4566]<=16'd0; ROM3[4566]<=16'd23770; ROM4[4566]<=16'd57276;
ROM1[4567]<=16'd4862; ROM2[4567]<=16'd0; ROM3[4567]<=16'd23769; ROM4[4567]<=16'd57272;
ROM1[4568]<=16'd4839; ROM2[4568]<=16'd0; ROM3[4568]<=16'd23768; ROM4[4568]<=16'd57269;
ROM1[4569]<=16'd4827; ROM2[4569]<=16'd0; ROM3[4569]<=16'd23776; ROM4[4569]<=16'd57275;
ROM1[4570]<=16'd4805; ROM2[4570]<=16'd0; ROM3[4570]<=16'd23778; ROM4[4570]<=16'd57269;
ROM1[4571]<=16'd4782; ROM2[4571]<=16'd0; ROM3[4571]<=16'd23766; ROM4[4571]<=16'd57253;
ROM1[4572]<=16'd4790; ROM2[4572]<=16'd0; ROM3[4572]<=16'd23769; ROM4[4572]<=16'd57258;
ROM1[4573]<=16'd4813; ROM2[4573]<=16'd0; ROM3[4573]<=16'd23759; ROM4[4573]<=16'd57259;
ROM1[4574]<=16'd4833; ROM2[4574]<=16'd0; ROM3[4574]<=16'd23736; ROM4[4574]<=16'd57246;
ROM1[4575]<=16'd4838; ROM2[4575]<=16'd0; ROM3[4575]<=16'd23741; ROM4[4575]<=16'd57253;
ROM1[4576]<=16'd4821; ROM2[4576]<=16'd0; ROM3[4576]<=16'd23749; ROM4[4576]<=16'd57252;
ROM1[4577]<=16'd4796; ROM2[4577]<=16'd0; ROM3[4577]<=16'd23750; ROM4[4577]<=16'd57241;
ROM1[4578]<=16'd4786; ROM2[4578]<=16'd0; ROM3[4578]<=16'd23765; ROM4[4578]<=16'd57249;
ROM1[4579]<=16'd4777; ROM2[4579]<=16'd0; ROM3[4579]<=16'd23778; ROM4[4579]<=16'd57257;
ROM1[4580]<=16'd4771; ROM2[4580]<=16'd0; ROM3[4580]<=16'd23765; ROM4[4580]<=16'd57247;
ROM1[4581]<=16'd4790; ROM2[4581]<=16'd0; ROM3[4581]<=16'd23754; ROM4[4581]<=16'd57241;
ROM1[4582]<=16'd4817; ROM2[4582]<=16'd0; ROM3[4582]<=16'd23738; ROM4[4582]<=16'd57234;
ROM1[4583]<=16'd4823; ROM2[4583]<=16'd0; ROM3[4583]<=16'd23727; ROM4[4583]<=16'd57231;
ROM1[4584]<=16'd4818; ROM2[4584]<=16'd0; ROM3[4584]<=16'd23736; ROM4[4584]<=16'd57238;
ROM1[4585]<=16'd4806; ROM2[4585]<=16'd0; ROM3[4585]<=16'd23747; ROM4[4585]<=16'd57243;
ROM1[4586]<=16'd4795; ROM2[4586]<=16'd0; ROM3[4586]<=16'd23752; ROM4[4586]<=16'd57242;
ROM1[4587]<=16'd4771; ROM2[4587]<=16'd0; ROM3[4587]<=16'd23746; ROM4[4587]<=16'd57232;
ROM1[4588]<=16'd4768; ROM2[4588]<=16'd0; ROM3[4588]<=16'd23746; ROM4[4588]<=16'd57227;
ROM1[4589]<=16'd4800; ROM2[4589]<=16'd0; ROM3[4589]<=16'd23751; ROM4[4589]<=16'd57241;
ROM1[4590]<=16'd4828; ROM2[4590]<=16'd0; ROM3[4590]<=16'd23734; ROM4[4590]<=16'd57240;
ROM1[4591]<=16'd4828; ROM2[4591]<=16'd0; ROM3[4591]<=16'd23709; ROM4[4591]<=16'd57226;
ROM1[4592]<=16'd4817; ROM2[4592]<=16'd0; ROM3[4592]<=16'd23715; ROM4[4592]<=16'd57229;
ROM1[4593]<=16'd4795; ROM2[4593]<=16'd0; ROM3[4593]<=16'd23714; ROM4[4593]<=16'd57222;
ROM1[4594]<=16'd4784; ROM2[4594]<=16'd0; ROM3[4594]<=16'd23725; ROM4[4594]<=16'd57223;
ROM1[4595]<=16'd4784; ROM2[4595]<=16'd0; ROM3[4595]<=16'd23748; ROM4[4595]<=16'd57235;
ROM1[4596]<=16'd4784; ROM2[4596]<=16'd0; ROM3[4596]<=16'd23758; ROM4[4596]<=16'd57243;
ROM1[4597]<=16'd4785; ROM2[4597]<=16'd0; ROM3[4597]<=16'd23752; ROM4[4597]<=16'd57240;
ROM1[4598]<=16'd4810; ROM2[4598]<=16'd0; ROM3[4598]<=16'd23741; ROM4[4598]<=16'd57242;
ROM1[4599]<=16'd4851; ROM2[4599]<=16'd0; ROM3[4599]<=16'd23745; ROM4[4599]<=16'd57258;
ROM1[4600]<=16'd4852; ROM2[4600]<=16'd0; ROM3[4600]<=16'd23747; ROM4[4600]<=16'd57262;
ROM1[4601]<=16'd4835; ROM2[4601]<=16'd0; ROM3[4601]<=16'd23751; ROM4[4601]<=16'd57261;
ROM1[4602]<=16'd4812; ROM2[4602]<=16'd0; ROM3[4602]<=16'd23754; ROM4[4602]<=16'd57253;
ROM1[4603]<=16'd4799; ROM2[4603]<=16'd0; ROM3[4603]<=16'd23753; ROM4[4603]<=16'd57249;
ROM1[4604]<=16'd4776; ROM2[4604]<=16'd0; ROM3[4604]<=16'd23743; ROM4[4604]<=16'd57238;
ROM1[4605]<=16'd4766; ROM2[4605]<=16'd0; ROM3[4605]<=16'd23730; ROM4[4605]<=16'd57227;
ROM1[4606]<=16'd4785; ROM2[4606]<=16'd0; ROM3[4606]<=16'd23723; ROM4[4606]<=16'd57223;
ROM1[4607]<=16'd4812; ROM2[4607]<=16'd0; ROM3[4607]<=16'd23711; ROM4[4607]<=16'd57218;
ROM1[4608]<=16'd4822; ROM2[4608]<=16'd0; ROM3[4608]<=16'd23715; ROM4[4608]<=16'd57224;
ROM1[4609]<=16'd4821; ROM2[4609]<=16'd0; ROM3[4609]<=16'd23732; ROM4[4609]<=16'd57239;
ROM1[4610]<=16'd4802; ROM2[4610]<=16'd0; ROM3[4610]<=16'd23739; ROM4[4610]<=16'd57240;
ROM1[4611]<=16'd4763; ROM2[4611]<=16'd0; ROM3[4611]<=16'd23724; ROM4[4611]<=16'd57215;
ROM1[4612]<=16'd4738; ROM2[4612]<=16'd0; ROM3[4612]<=16'd23716; ROM4[4612]<=16'd57199;
ROM1[4613]<=16'd4740; ROM2[4613]<=16'd0; ROM3[4613]<=16'd23725; ROM4[4613]<=16'd57205;
ROM1[4614]<=16'd4767; ROM2[4614]<=16'd0; ROM3[4614]<=16'd23736; ROM4[4614]<=16'd57220;
ROM1[4615]<=16'd4805; ROM2[4615]<=16'd0; ROM3[4615]<=16'd23730; ROM4[4615]<=16'd57227;
ROM1[4616]<=16'd4821; ROM2[4616]<=16'd0; ROM3[4616]<=16'd23723; ROM4[4616]<=16'd57225;
ROM1[4617]<=16'd4806; ROM2[4617]<=16'd0; ROM3[4617]<=16'd23716; ROM4[4617]<=16'd57219;
ROM1[4618]<=16'd4789; ROM2[4618]<=16'd0; ROM3[4618]<=16'd23717; ROM4[4618]<=16'd57219;
ROM1[4619]<=16'd4793; ROM2[4619]<=16'd0; ROM3[4619]<=16'd23745; ROM4[4619]<=16'd57240;
ROM1[4620]<=16'd4806; ROM2[4620]<=16'd0; ROM3[4620]<=16'd23775; ROM4[4620]<=16'd57263;
ROM1[4621]<=16'd4775; ROM2[4621]<=16'd0; ROM3[4621]<=16'd23761; ROM4[4621]<=16'd57243;
ROM1[4622]<=16'd4765; ROM2[4622]<=16'd0; ROM3[4622]<=16'd23734; ROM4[4622]<=16'd57225;
ROM1[4623]<=16'd4803; ROM2[4623]<=16'd0; ROM3[4623]<=16'd23728; ROM4[4623]<=16'd57236;
ROM1[4624]<=16'd4836; ROM2[4624]<=16'd0; ROM3[4624]<=16'd23725; ROM4[4624]<=16'd57246;
ROM1[4625]<=16'd4849; ROM2[4625]<=16'd0; ROM3[4625]<=16'd23740; ROM4[4625]<=16'd57264;
ROM1[4626]<=16'd4840; ROM2[4626]<=16'd0; ROM3[4626]<=16'd23757; ROM4[4626]<=16'd57272;
ROM1[4627]<=16'd4819; ROM2[4627]<=16'd0; ROM3[4627]<=16'd23767; ROM4[4627]<=16'd57271;
ROM1[4628]<=16'd4802; ROM2[4628]<=16'd0; ROM3[4628]<=16'd23766; ROM4[4628]<=16'd57269;
ROM1[4629]<=16'd4795; ROM2[4629]<=16'd0; ROM3[4629]<=16'd23780; ROM4[4629]<=16'd57272;
ROM1[4630]<=16'd4810; ROM2[4630]<=16'd0; ROM3[4630]<=16'd23797; ROM4[4630]<=16'd57284;
ROM1[4631]<=16'd4824; ROM2[4631]<=16'd0; ROM3[4631]<=16'd23782; ROM4[4631]<=16'd57275;
ROM1[4632]<=16'd4842; ROM2[4632]<=16'd0; ROM3[4632]<=16'd23761; ROM4[4632]<=16'd57258;
ROM1[4633]<=16'd4852; ROM2[4633]<=16'd0; ROM3[4633]<=16'd23759; ROM4[4633]<=16'd57258;
ROM1[4634]<=16'd4851; ROM2[4634]<=16'd0; ROM3[4634]<=16'd23778; ROM4[4634]<=16'd57275;
ROM1[4635]<=16'd4849; ROM2[4635]<=16'd0; ROM3[4635]<=16'd23803; ROM4[4635]<=16'd57295;
ROM1[4636]<=16'd4820; ROM2[4636]<=16'd0; ROM3[4636]<=16'd23791; ROM4[4636]<=16'd57281;
ROM1[4637]<=16'd4778; ROM2[4637]<=16'd0; ROM3[4637]<=16'd23769; ROM4[4637]<=16'd57254;
ROM1[4638]<=16'd4766; ROM2[4638]<=16'd0; ROM3[4638]<=16'd23759; ROM4[4638]<=16'd57247;
ROM1[4639]<=16'd4784; ROM2[4639]<=16'd0; ROM3[4639]<=16'd23752; ROM4[4639]<=16'd57246;
ROM1[4640]<=16'd4831; ROM2[4640]<=16'd0; ROM3[4640]<=16'd23755; ROM4[4640]<=16'd57262;
ROM1[4641]<=16'd4859; ROM2[4641]<=16'd0; ROM3[4641]<=16'd23756; ROM4[4641]<=16'd57273;
ROM1[4642]<=16'd4839; ROM2[4642]<=16'd0; ROM3[4642]<=16'd23749; ROM4[4642]<=16'd57264;
ROM1[4643]<=16'd4815; ROM2[4643]<=16'd0; ROM3[4643]<=16'd23754; ROM4[4643]<=16'd57257;
ROM1[4644]<=16'd4805; ROM2[4644]<=16'd0; ROM3[4644]<=16'd23767; ROM4[4644]<=16'd57262;
ROM1[4645]<=16'd4795; ROM2[4645]<=16'd0; ROM3[4645]<=16'd23777; ROM4[4645]<=16'd57267;
ROM1[4646]<=16'd4780; ROM2[4646]<=16'd0; ROM3[4646]<=16'd23779; ROM4[4646]<=16'd57261;
ROM1[4647]<=16'd4787; ROM2[4647]<=16'd0; ROM3[4647]<=16'd23777; ROM4[4647]<=16'd57263;
ROM1[4648]<=16'd4823; ROM2[4648]<=16'd0; ROM3[4648]<=16'd23778; ROM4[4648]<=16'd57271;
ROM1[4649]<=16'd4848; ROM2[4649]<=16'd0; ROM3[4649]<=16'd23767; ROM4[4649]<=16'd57274;
ROM1[4650]<=16'd4841; ROM2[4650]<=16'd0; ROM3[4650]<=16'd23758; ROM4[4650]<=16'd57268;
ROM1[4651]<=16'd4824; ROM2[4651]<=16'd0; ROM3[4651]<=16'd23762; ROM4[4651]<=16'd57265;
ROM1[4652]<=16'd4802; ROM2[4652]<=16'd0; ROM3[4652]<=16'd23765; ROM4[4652]<=16'd57259;
ROM1[4653]<=16'd4783; ROM2[4653]<=16'd0; ROM3[4653]<=16'd23763; ROM4[4653]<=16'd57251;
ROM1[4654]<=16'd4775; ROM2[4654]<=16'd0; ROM3[4654]<=16'd23766; ROM4[4654]<=16'd57255;
ROM1[4655]<=16'd4775; ROM2[4655]<=16'd0; ROM3[4655]<=16'd23759; ROM4[4655]<=16'd57252;
ROM1[4656]<=16'd4794; ROM2[4656]<=16'd0; ROM3[4656]<=16'd23741; ROM4[4656]<=16'd57241;
ROM1[4657]<=16'd4834; ROM2[4657]<=16'd0; ROM3[4657]<=16'd23726; ROM4[4657]<=16'd57242;
ROM1[4658]<=16'd4846; ROM2[4658]<=16'd0; ROM3[4658]<=16'd23722; ROM4[4658]<=16'd57243;
ROM1[4659]<=16'd4837; ROM2[4659]<=16'd0; ROM3[4659]<=16'd23734; ROM4[4659]<=16'd57244;
ROM1[4660]<=16'd4816; ROM2[4660]<=16'd0; ROM3[4660]<=16'd23744; ROM4[4660]<=16'd57246;
ROM1[4661]<=16'd4803; ROM2[4661]<=16'd0; ROM3[4661]<=16'd23750; ROM4[4661]<=16'd57245;
ROM1[4662]<=16'd4793; ROM2[4662]<=16'd0; ROM3[4662]<=16'd23758; ROM4[4662]<=16'd57248;
ROM1[4663]<=16'd4785; ROM2[4663]<=16'd0; ROM3[4663]<=16'd23761; ROM4[4663]<=16'd57247;
ROM1[4664]<=16'd4798; ROM2[4664]<=16'd0; ROM3[4664]<=16'd23749; ROM4[4664]<=16'd57244;
ROM1[4665]<=16'd4825; ROM2[4665]<=16'd0; ROM3[4665]<=16'd23733; ROM4[4665]<=16'd57239;
ROM1[4666]<=16'd4846; ROM2[4666]<=16'd0; ROM3[4666]<=16'd23735; ROM4[4666]<=16'd57247;
ROM1[4667]<=16'd4860; ROM2[4667]<=16'd0; ROM3[4667]<=16'd23753; ROM4[4667]<=16'd57270;
ROM1[4668]<=16'd4854; ROM2[4668]<=16'd0; ROM3[4668]<=16'd23770; ROM4[4668]<=16'd57279;
ROM1[4669]<=16'd4825; ROM2[4669]<=16'd0; ROM3[4669]<=16'd23770; ROM4[4669]<=16'd57272;
ROM1[4670]<=16'd4810; ROM2[4670]<=16'd0; ROM3[4670]<=16'd23772; ROM4[4670]<=16'd57271;
ROM1[4671]<=16'd4790; ROM2[4671]<=16'd0; ROM3[4671]<=16'd23758; ROM4[4671]<=16'd57256;
ROM1[4672]<=16'd4782; ROM2[4672]<=16'd0; ROM3[4672]<=16'd23737; ROM4[4672]<=16'd57242;
ROM1[4673]<=16'd4824; ROM2[4673]<=16'd0; ROM3[4673]<=16'd23738; ROM4[4673]<=16'd57258;
ROM1[4674]<=16'd4849; ROM2[4674]<=16'd0; ROM3[4674]<=16'd23728; ROM4[4674]<=16'd57259;
ROM1[4675]<=16'd4850; ROM2[4675]<=16'd0; ROM3[4675]<=16'd23733; ROM4[4675]<=16'd57263;
ROM1[4676]<=16'd4856; ROM2[4676]<=16'd0; ROM3[4676]<=16'd23759; ROM4[4676]<=16'd57281;
ROM1[4677]<=16'd4839; ROM2[4677]<=16'd0; ROM3[4677]<=16'd23774; ROM4[4677]<=16'd57284;
ROM1[4678]<=16'd4820; ROM2[4678]<=16'd0; ROM3[4678]<=16'd23778; ROM4[4678]<=16'd57280;
ROM1[4679]<=16'd4800; ROM2[4679]<=16'd0; ROM3[4679]<=16'd23775; ROM4[4679]<=16'd57273;
ROM1[4680]<=16'd4795; ROM2[4680]<=16'd0; ROM3[4680]<=16'd23773; ROM4[4680]<=16'd57269;
ROM1[4681]<=16'd4826; ROM2[4681]<=16'd0; ROM3[4681]<=16'd23773; ROM4[4681]<=16'd57274;
ROM1[4682]<=16'd4866; ROM2[4682]<=16'd0; ROM3[4682]<=16'd23769; ROM4[4682]<=16'd57282;
ROM1[4683]<=16'd4878; ROM2[4683]<=16'd0; ROM3[4683]<=16'd23770; ROM4[4683]<=16'd57283;
ROM1[4684]<=16'd4857; ROM2[4684]<=16'd0; ROM3[4684]<=16'd23766; ROM4[4684]<=16'd57277;
ROM1[4685]<=16'd4833; ROM2[4685]<=16'd0; ROM3[4685]<=16'd23769; ROM4[4685]<=16'd57277;
ROM1[4686]<=16'd4825; ROM2[4686]<=16'd0; ROM3[4686]<=16'd23782; ROM4[4686]<=16'd57280;
ROM1[4687]<=16'd4814; ROM2[4687]<=16'd0; ROM3[4687]<=16'd23794; ROM4[4687]<=16'd57287;
ROM1[4688]<=16'd4823; ROM2[4688]<=16'd0; ROM3[4688]<=16'd23806; ROM4[4688]<=16'd57301;
ROM1[4689]<=16'd4858; ROM2[4689]<=16'd0; ROM3[4689]<=16'd23816; ROM4[4689]<=16'd57314;
ROM1[4690]<=16'd4896; ROM2[4690]<=16'd0; ROM3[4690]<=16'd23804; ROM4[4690]<=16'd57314;
ROM1[4691]<=16'd4918; ROM2[4691]<=16'd0; ROM3[4691]<=16'd23795; ROM4[4691]<=16'd57316;
ROM1[4692]<=16'd4901; ROM2[4692]<=16'd0; ROM3[4692]<=16'd23790; ROM4[4692]<=16'd57309;
ROM1[4693]<=16'd4859; ROM2[4693]<=16'd0; ROM3[4693]<=16'd23776; ROM4[4693]<=16'd57291;
ROM1[4694]<=16'd4843; ROM2[4694]<=16'd0; ROM3[4694]<=16'd23783; ROM4[4694]<=16'd57292;
ROM1[4695]<=16'd4837; ROM2[4695]<=16'd0; ROM3[4695]<=16'd23797; ROM4[4695]<=16'd57298;
ROM1[4696]<=16'd4841; ROM2[4696]<=16'd0; ROM3[4696]<=16'd23806; ROM4[4696]<=16'd57306;
ROM1[4697]<=16'd4858; ROM2[4697]<=16'd0; ROM3[4697]<=16'd23804; ROM4[4697]<=16'd57308;
ROM1[4698]<=16'd4880; ROM2[4698]<=16'd0; ROM3[4698]<=16'd23788; ROM4[4698]<=16'd57300;
ROM1[4699]<=16'd4901; ROM2[4699]<=16'd0; ROM3[4699]<=16'd23774; ROM4[4699]<=16'd57297;
ROM1[4700]<=16'd4902; ROM2[4700]<=16'd0; ROM3[4700]<=16'd23779; ROM4[4700]<=16'd57303;
ROM1[4701]<=16'd4888; ROM2[4701]<=16'd0; ROM3[4701]<=16'd23791; ROM4[4701]<=16'd57306;
ROM1[4702]<=16'd4872; ROM2[4702]<=16'd0; ROM3[4702]<=16'd23801; ROM4[4702]<=16'd57307;
ROM1[4703]<=16'd4858; ROM2[4703]<=16'd0; ROM3[4703]<=16'd23810; ROM4[4703]<=16'd57310;
ROM1[4704]<=16'd4842; ROM2[4704]<=16'd0; ROM3[4704]<=16'd23817; ROM4[4704]<=16'd57308;
ROM1[4705]<=16'd4838; ROM2[4705]<=16'd0; ROM3[4705]<=16'd23815; ROM4[4705]<=16'd57302;
ROM1[4706]<=16'd4852; ROM2[4706]<=16'd0; ROM3[4706]<=16'd23802; ROM4[4706]<=16'd57297;
ROM1[4707]<=16'd4874; ROM2[4707]<=16'd0; ROM3[4707]<=16'd23784; ROM4[4707]<=16'd57290;
ROM1[4708]<=16'd4879; ROM2[4708]<=16'd0; ROM3[4708]<=16'd23782; ROM4[4708]<=16'd57291;
ROM1[4709]<=16'd4871; ROM2[4709]<=16'd0; ROM3[4709]<=16'd23792; ROM4[4709]<=16'd57294;
ROM1[4710]<=16'd4853; ROM2[4710]<=16'd0; ROM3[4710]<=16'd23802; ROM4[4710]<=16'd57296;
ROM1[4711]<=16'd4851; ROM2[4711]<=16'd0; ROM3[4711]<=16'd23821; ROM4[4711]<=16'd57305;
ROM1[4712]<=16'd4852; ROM2[4712]<=16'd0; ROM3[4712]<=16'd23842; ROM4[4712]<=16'd57321;
ROM1[4713]<=16'd4828; ROM2[4713]<=16'd0; ROM3[4713]<=16'd23828; ROM4[4713]<=16'd57305;
ROM1[4714]<=16'd4824; ROM2[4714]<=16'd0; ROM3[4714]<=16'd23805; ROM4[4714]<=16'd57289;
ROM1[4715]<=16'd4857; ROM2[4715]<=16'd0; ROM3[4715]<=16'd23794; ROM4[4715]<=16'd57289;
ROM1[4716]<=16'd4878; ROM2[4716]<=16'd0; ROM3[4716]<=16'd23787; ROM4[4716]<=16'd57291;
ROM1[4717]<=16'd4894; ROM2[4717]<=16'd0; ROM3[4717]<=16'd23811; ROM4[4717]<=16'd57313;
ROM1[4718]<=16'd4899; ROM2[4718]<=16'd0; ROM3[4718]<=16'd23839; ROM4[4718]<=16'd57332;
ROM1[4719]<=16'd4868; ROM2[4719]<=16'd0; ROM3[4719]<=16'd23827; ROM4[4719]<=16'd57316;
ROM1[4720]<=16'd4833; ROM2[4720]<=16'd0; ROM3[4720]<=16'd23811; ROM4[4720]<=16'd57295;
ROM1[4721]<=16'd4831; ROM2[4721]<=16'd0; ROM3[4721]<=16'd23816; ROM4[4721]<=16'd57300;
ROM1[4722]<=16'd4841; ROM2[4722]<=16'd0; ROM3[4722]<=16'd23811; ROM4[4722]<=16'd57305;
ROM1[4723]<=16'd4864; ROM2[4723]<=16'd0; ROM3[4723]<=16'd23798; ROM4[4723]<=16'd57303;
ROM1[4724]<=16'd4889; ROM2[4724]<=16'd0; ROM3[4724]<=16'd23779; ROM4[4724]<=16'd57297;
ROM1[4725]<=16'd4879; ROM2[4725]<=16'd0; ROM3[4725]<=16'd23779; ROM4[4725]<=16'd57301;
ROM1[4726]<=16'd4870; ROM2[4726]<=16'd0; ROM3[4726]<=16'd23795; ROM4[4726]<=16'd57311;
ROM1[4727]<=16'd4863; ROM2[4727]<=16'd0; ROM3[4727]<=16'd23812; ROM4[4727]<=16'd57318;
ROM1[4728]<=16'd4840; ROM2[4728]<=16'd0; ROM3[4728]<=16'd23812; ROM4[4728]<=16'd57313;
ROM1[4729]<=16'd4829; ROM2[4729]<=16'd0; ROM3[4729]<=16'd23806; ROM4[4729]<=16'd57302;
ROM1[4730]<=16'd4840; ROM2[4730]<=16'd0; ROM3[4730]<=16'd23804; ROM4[4730]<=16'd57297;
ROM1[4731]<=16'd4874; ROM2[4731]<=16'd0; ROM3[4731]<=16'd23806; ROM4[4731]<=16'd57307;
ROM1[4732]<=16'd4902; ROM2[4732]<=16'd0; ROM3[4732]<=16'd23799; ROM4[4732]<=16'd57310;
ROM1[4733]<=16'd4899; ROM2[4733]<=16'd0; ROM3[4733]<=16'd23796; ROM4[4733]<=16'd57307;
ROM1[4734]<=16'd4880; ROM2[4734]<=16'd0; ROM3[4734]<=16'd23802; ROM4[4734]<=16'd57304;
ROM1[4735]<=16'd4853; ROM2[4735]<=16'd0; ROM3[4735]<=16'd23800; ROM4[4735]<=16'd57299;
ROM1[4736]<=16'd4859; ROM2[4736]<=16'd0; ROM3[4736]<=16'd23822; ROM4[4736]<=16'd57317;
ROM1[4737]<=16'd4865; ROM2[4737]<=16'd0; ROM3[4737]<=16'd23846; ROM4[4737]<=16'd57336;
ROM1[4738]<=16'd4852; ROM2[4738]<=16'd0; ROM3[4738]<=16'd23836; ROM4[4738]<=16'd57326;
ROM1[4739]<=16'd4850; ROM2[4739]<=16'd0; ROM3[4739]<=16'd23813; ROM4[4739]<=16'd57307;
ROM1[4740]<=16'd4882; ROM2[4740]<=16'd0; ROM3[4740]<=16'd23792; ROM4[4740]<=16'd57302;
ROM1[4741]<=16'd4902; ROM2[4741]<=16'd0; ROM3[4741]<=16'd23781; ROM4[4741]<=16'd57302;
ROM1[4742]<=16'd4896; ROM2[4742]<=16'd0; ROM3[4742]<=16'd23788; ROM4[4742]<=16'd57308;
ROM1[4743]<=16'd4888; ROM2[4743]<=16'd0; ROM3[4743]<=16'd23809; ROM4[4743]<=16'd57320;
ROM1[4744]<=16'd4870; ROM2[4744]<=16'd0; ROM3[4744]<=16'd23821; ROM4[4744]<=16'd57319;
ROM1[4745]<=16'd4841; ROM2[4745]<=16'd0; ROM3[4745]<=16'd23818; ROM4[4745]<=16'd57312;
ROM1[4746]<=16'd4826; ROM2[4746]<=16'd0; ROM3[4746]<=16'd23816; ROM4[4746]<=16'd57306;
ROM1[4747]<=16'd4834; ROM2[4747]<=16'd0; ROM3[4747]<=16'd23808; ROM4[4747]<=16'd57301;
ROM1[4748]<=16'd4862; ROM2[4748]<=16'd0; ROM3[4748]<=16'd23795; ROM4[4748]<=16'd57299;
ROM1[4749]<=16'd4884; ROM2[4749]<=16'd0; ROM3[4749]<=16'd23776; ROM4[4749]<=16'd57291;
ROM1[4750]<=16'd4868; ROM2[4750]<=16'd0; ROM3[4750]<=16'd23763; ROM4[4750]<=16'd57277;
ROM1[4751]<=16'd4849; ROM2[4751]<=16'd0; ROM3[4751]<=16'd23768; ROM4[4751]<=16'd57279;
ROM1[4752]<=16'd4843; ROM2[4752]<=16'd0; ROM3[4752]<=16'd23778; ROM4[4752]<=16'd57284;
ROM1[4753]<=16'd4838; ROM2[4753]<=16'd0; ROM3[4753]<=16'd23790; ROM4[4753]<=16'd57288;
ROM1[4754]<=16'd4830; ROM2[4754]<=16'd0; ROM3[4754]<=16'd23799; ROM4[4754]<=16'd57294;
ROM1[4755]<=16'd4814; ROM2[4755]<=16'd0; ROM3[4755]<=16'd23781; ROM4[4755]<=16'd57275;
ROM1[4756]<=16'd4810; ROM2[4756]<=16'd0; ROM3[4756]<=16'd23753; ROM4[4756]<=16'd57249;
ROM1[4757]<=16'd4834; ROM2[4757]<=16'd0; ROM3[4757]<=16'd23734; ROM4[4757]<=16'd57243;
ROM1[4758]<=16'd4842; ROM2[4758]<=16'd0; ROM3[4758]<=16'd23732; ROM4[4758]<=16'd57245;
ROM1[4759]<=16'd4836; ROM2[4759]<=16'd0; ROM3[4759]<=16'd23742; ROM4[4759]<=16'd57254;
ROM1[4760]<=16'd4828; ROM2[4760]<=16'd0; ROM3[4760]<=16'd23759; ROM4[4760]<=16'd57264;
ROM1[4761]<=16'd4817; ROM2[4761]<=16'd0; ROM3[4761]<=16'd23767; ROM4[4761]<=16'd57265;
ROM1[4762]<=16'd4802; ROM2[4762]<=16'd0; ROM3[4762]<=16'd23773; ROM4[4762]<=16'd57265;
ROM1[4763]<=16'd4810; ROM2[4763]<=16'd0; ROM3[4763]<=16'd23789; ROM4[4763]<=16'd57275;
ROM1[4764]<=16'd4827; ROM2[4764]<=16'd0; ROM3[4764]<=16'd23786; ROM4[4764]<=16'd57278;
ROM1[4765]<=16'd4864; ROM2[4765]<=16'd0; ROM3[4765]<=16'd23779; ROM4[4765]<=16'd57286;
ROM1[4766]<=16'd4890; ROM2[4766]<=16'd0; ROM3[4766]<=16'd23779; ROM4[4766]<=16'd57295;
ROM1[4767]<=16'd4879; ROM2[4767]<=16'd0; ROM3[4767]<=16'd23782; ROM4[4767]<=16'd57295;
ROM1[4768]<=16'd4862; ROM2[4768]<=16'd0; ROM3[4768]<=16'd23792; ROM4[4768]<=16'd57295;
ROM1[4769]<=16'd4844; ROM2[4769]<=16'd0; ROM3[4769]<=16'd23797; ROM4[4769]<=16'd57291;
ROM1[4770]<=16'd4826; ROM2[4770]<=16'd0; ROM3[4770]<=16'd23801; ROM4[4770]<=16'd57288;
ROM1[4771]<=16'd4826; ROM2[4771]<=16'd0; ROM3[4771]<=16'd23809; ROM4[4771]<=16'd57291;
ROM1[4772]<=16'd4859; ROM2[4772]<=16'd0; ROM3[4772]<=16'd23822; ROM4[4772]<=16'd57313;
ROM1[4773]<=16'd4890; ROM2[4773]<=16'd0; ROM3[4773]<=16'd23815; ROM4[4773]<=16'd57321;
ROM1[4774]<=16'd4898; ROM2[4774]<=16'd0; ROM3[4774]<=16'd23788; ROM4[4774]<=16'd57305;
ROM1[4775]<=16'd4878; ROM2[4775]<=16'd0; ROM3[4775]<=16'd23773; ROM4[4775]<=16'd57292;
ROM1[4776]<=16'd4854; ROM2[4776]<=16'd0; ROM3[4776]<=16'd23777; ROM4[4776]<=16'd57283;
ROM1[4777]<=16'd4845; ROM2[4777]<=16'd0; ROM3[4777]<=16'd23789; ROM4[4777]<=16'd57281;
ROM1[4778]<=16'd4842; ROM2[4778]<=16'd0; ROM3[4778]<=16'd23797; ROM4[4778]<=16'd57288;
ROM1[4779]<=16'd4830; ROM2[4779]<=16'd0; ROM3[4779]<=16'd23802; ROM4[4779]<=16'd57289;
ROM1[4780]<=16'd4826; ROM2[4780]<=16'd0; ROM3[4780]<=16'd23795; ROM4[4780]<=16'd57284;
ROM1[4781]<=16'd4841; ROM2[4781]<=16'd0; ROM3[4781]<=16'd23778; ROM4[4781]<=16'd57279;
ROM1[4782]<=16'd4875; ROM2[4782]<=16'd0; ROM3[4782]<=16'd23771; ROM4[4782]<=16'd57282;
ROM1[4783]<=16'd4886; ROM2[4783]<=16'd0; ROM3[4783]<=16'd23775; ROM4[4783]<=16'd57286;
ROM1[4784]<=16'd4870; ROM2[4784]<=16'd0; ROM3[4784]<=16'd23778; ROM4[4784]<=16'd57285;
ROM1[4785]<=16'd4851; ROM2[4785]<=16'd0; ROM3[4785]<=16'd23792; ROM4[4785]<=16'd57288;
ROM1[4786]<=16'd4843; ROM2[4786]<=16'd0; ROM3[4786]<=16'd23808; ROM4[4786]<=16'd57294;
ROM1[4787]<=16'd4834; ROM2[4787]<=16'd0; ROM3[4787]<=16'd23816; ROM4[4787]<=16'd57299;
ROM1[4788]<=16'd4836; ROM2[4788]<=16'd0; ROM3[4788]<=16'd23818; ROM4[4788]<=16'd57300;
ROM1[4789]<=16'd4852; ROM2[4789]<=16'd0; ROM3[4789]<=16'd23810; ROM4[4789]<=16'd57299;
ROM1[4790]<=16'd4889; ROM2[4790]<=16'd0; ROM3[4790]<=16'd23804; ROM4[4790]<=16'd57302;
ROM1[4791]<=16'd4908; ROM2[4791]<=16'd0; ROM3[4791]<=16'd23794; ROM4[4791]<=16'd57296;
ROM1[4792]<=16'd4888; ROM2[4792]<=16'd0; ROM3[4792]<=16'd23788; ROM4[4792]<=16'd57290;
ROM1[4793]<=16'd4891; ROM2[4793]<=16'd0; ROM3[4793]<=16'd23817; ROM4[4793]<=16'd57313;
ROM1[4794]<=16'd4890; ROM2[4794]<=16'd0; ROM3[4794]<=16'd23833; ROM4[4794]<=16'd57322;
ROM1[4795]<=16'd4849; ROM2[4795]<=16'd0; ROM3[4795]<=16'd23809; ROM4[4795]<=16'd57296;
ROM1[4796]<=16'd4814; ROM2[4796]<=16'd0; ROM3[4796]<=16'd23785; ROM4[4796]<=16'd57271;
ROM1[4797]<=16'd4814; ROM2[4797]<=16'd0; ROM3[4797]<=16'd23774; ROM4[4797]<=16'd57261;
ROM1[4798]<=16'd4844; ROM2[4798]<=16'd0; ROM3[4798]<=16'd23770; ROM4[4798]<=16'd57265;
ROM1[4799]<=16'd4890; ROM2[4799]<=16'd0; ROM3[4799]<=16'd23778; ROM4[4799]<=16'd57288;
ROM1[4800]<=16'd4902; ROM2[4800]<=16'd0; ROM3[4800]<=16'd23794; ROM4[4800]<=16'd57304;
ROM1[4801]<=16'd4880; ROM2[4801]<=16'd0; ROM3[4801]<=16'd23798; ROM4[4801]<=16'd57298;
ROM1[4802]<=16'd4864; ROM2[4802]<=16'd0; ROM3[4802]<=16'd23804; ROM4[4802]<=16'd57300;
ROM1[4803]<=16'd4859; ROM2[4803]<=16'd0; ROM3[4803]<=16'd23820; ROM4[4803]<=16'd57313;
ROM1[4804]<=16'd4851; ROM2[4804]<=16'd0; ROM3[4804]<=16'd23831; ROM4[4804]<=16'd57318;
ROM1[4805]<=16'd4849; ROM2[4805]<=16'd0; ROM3[4805]<=16'd23825; ROM4[4805]<=16'd57310;
ROM1[4806]<=16'd4857; ROM2[4806]<=16'd0; ROM3[4806]<=16'd23798; ROM4[4806]<=16'd57292;
ROM1[4807]<=16'd4880; ROM2[4807]<=16'd0; ROM3[4807]<=16'd23776; ROM4[4807]<=16'd57285;
ROM1[4808]<=16'd4894; ROM2[4808]<=16'd0; ROM3[4808]<=16'd23780; ROM4[4808]<=16'd57292;
ROM1[4809]<=16'd4890; ROM2[4809]<=16'd0; ROM3[4809]<=16'd23790; ROM4[4809]<=16'd57303;
ROM1[4810]<=16'd4885; ROM2[4810]<=16'd0; ROM3[4810]<=16'd23812; ROM4[4810]<=16'd57318;
ROM1[4811]<=16'd4886; ROM2[4811]<=16'd0; ROM3[4811]<=16'd23834; ROM4[4811]<=16'd57331;
ROM1[4812]<=16'd4860; ROM2[4812]<=16'd0; ROM3[4812]<=16'd23826; ROM4[4812]<=16'd57318;
ROM1[4813]<=16'd4827; ROM2[4813]<=16'd0; ROM3[4813]<=16'd23804; ROM4[4813]<=16'd57289;
ROM1[4814]<=16'd4829; ROM2[4814]<=16'd0; ROM3[4814]<=16'd23787; ROM4[4814]<=16'd57278;
ROM1[4815]<=16'd4856; ROM2[4815]<=16'd0; ROM3[4815]<=16'd23771; ROM4[4815]<=16'd57272;
ROM1[4816]<=16'd4875; ROM2[4816]<=16'd0; ROM3[4816]<=16'd23767; ROM4[4816]<=16'd57276;
ROM1[4817]<=16'd4868; ROM2[4817]<=16'd0; ROM3[4817]<=16'd23771; ROM4[4817]<=16'd57283;
ROM1[4818]<=16'd4851; ROM2[4818]<=16'd0; ROM3[4818]<=16'd23781; ROM4[4818]<=16'd57287;
ROM1[4819]<=16'd4839; ROM2[4819]<=16'd0; ROM3[4819]<=16'd23793; ROM4[4819]<=16'd57290;
ROM1[4820]<=16'd4836; ROM2[4820]<=16'd0; ROM3[4820]<=16'd23814; ROM4[4820]<=16'd57301;
ROM1[4821]<=16'd4844; ROM2[4821]<=16'd0; ROM3[4821]<=16'd23835; ROM4[4821]<=16'd57318;
ROM1[4822]<=16'd4858; ROM2[4822]<=16'd0; ROM3[4822]<=16'd23836; ROM4[4822]<=16'd57322;
ROM1[4823]<=16'd4876; ROM2[4823]<=16'd0; ROM3[4823]<=16'd23821; ROM4[4823]<=16'd57311;
ROM1[4824]<=16'd4891; ROM2[4824]<=16'd0; ROM3[4824]<=16'd23801; ROM4[4824]<=16'd57300;
ROM1[4825]<=16'd4887; ROM2[4825]<=16'd0; ROM3[4825]<=16'd23798; ROM4[4825]<=16'd57300;
ROM1[4826]<=16'd4866; ROM2[4826]<=16'd0; ROM3[4826]<=16'd23802; ROM4[4826]<=16'd57296;
ROM1[4827]<=16'd4849; ROM2[4827]<=16'd0; ROM3[4827]<=16'd23808; ROM4[4827]<=16'd57294;
ROM1[4828]<=16'd4841; ROM2[4828]<=16'd0; ROM3[4828]<=16'd23819; ROM4[4828]<=16'd57301;
ROM1[4829]<=16'd4841; ROM2[4829]<=16'd0; ROM3[4829]<=16'd23839; ROM4[4829]<=16'd57310;
ROM1[4830]<=16'd4838; ROM2[4830]<=16'd0; ROM3[4830]<=16'd23827; ROM4[4830]<=16'd57302;
ROM1[4831]<=16'd4844; ROM2[4831]<=16'd0; ROM3[4831]<=16'd23803; ROM4[4831]<=16'd57286;
ROM1[4832]<=16'd4880; ROM2[4832]<=16'd0; ROM3[4832]<=16'd23797; ROM4[4832]<=16'd57291;
ROM1[4833]<=16'd4888; ROM2[4833]<=16'd0; ROM3[4833]<=16'd23792; ROM4[4833]<=16'd57295;
ROM1[4834]<=16'd4870; ROM2[4834]<=16'd0; ROM3[4834]<=16'd23802; ROM4[4834]<=16'd57296;
ROM1[4835]<=16'd4856; ROM2[4835]<=16'd0; ROM3[4835]<=16'd23816; ROM4[4835]<=16'd57300;
ROM1[4836]<=16'd4860; ROM2[4836]<=16'd0; ROM3[4836]<=16'd23830; ROM4[4836]<=16'd57308;
ROM1[4837]<=16'd4878; ROM2[4837]<=16'd0; ROM3[4837]<=16'd23866; ROM4[4837]<=16'd57338;
ROM1[4838]<=16'd4879; ROM2[4838]<=16'd0; ROM3[4838]<=16'd23868; ROM4[4838]<=16'd57337;
ROM1[4839]<=16'd4857; ROM2[4839]<=16'd0; ROM3[4839]<=16'd23826; ROM4[4839]<=16'd57300;
ROM1[4840]<=16'd4874; ROM2[4840]<=16'd0; ROM3[4840]<=16'd23804; ROM4[4840]<=16'd57290;
ROM1[4841]<=16'd4870; ROM2[4841]<=16'd0; ROM3[4841]<=16'd23775; ROM4[4841]<=16'd57271;
ROM1[4842]<=16'd4861; ROM2[4842]<=16'd0; ROM3[4842]<=16'd23778; ROM4[4842]<=16'd57275;
ROM1[4843]<=16'd4870; ROM2[4843]<=16'd0; ROM3[4843]<=16'd23814; ROM4[4843]<=16'd57306;
ROM1[4844]<=16'd4859; ROM2[4844]<=16'd0; ROM3[4844]<=16'd23828; ROM4[4844]<=16'd57311;
ROM1[4845]<=16'd4831; ROM2[4845]<=16'd0; ROM3[4845]<=16'd23817; ROM4[4845]<=16'd57294;
ROM1[4846]<=16'd4814; ROM2[4846]<=16'd0; ROM3[4846]<=16'd23812; ROM4[4846]<=16'd57287;
ROM1[4847]<=16'd4834; ROM2[4847]<=16'd0; ROM3[4847]<=16'd23819; ROM4[4847]<=16'd57298;
ROM1[4848]<=16'd4863; ROM2[4848]<=16'd0; ROM3[4848]<=16'd23804; ROM4[4848]<=16'd57296;
ROM1[4849]<=16'd4889; ROM2[4849]<=16'd0; ROM3[4849]<=16'd23791; ROM4[4849]<=16'd57294;
ROM1[4850]<=16'd4890; ROM2[4850]<=16'd0; ROM3[4850]<=16'd23793; ROM4[4850]<=16'd57302;
ROM1[4851]<=16'd4875; ROM2[4851]<=16'd0; ROM3[4851]<=16'd23804; ROM4[4851]<=16'd57307;
ROM1[4852]<=16'd4859; ROM2[4852]<=16'd0; ROM3[4852]<=16'd23814; ROM4[4852]<=16'd57310;
ROM1[4853]<=16'd4836; ROM2[4853]<=16'd0; ROM3[4853]<=16'd23812; ROM4[4853]<=16'd57302;
ROM1[4854]<=16'd4796; ROM2[4854]<=16'd0; ROM3[4854]<=16'd23796; ROM4[4854]<=16'd57279;
ROM1[4855]<=16'd4798; ROM2[4855]<=16'd0; ROM3[4855]<=16'd23786; ROM4[4855]<=16'd57270;
ROM1[4856]<=16'd4821; ROM2[4856]<=16'd0; ROM3[4856]<=16'd23776; ROM4[4856]<=16'd57268;
ROM1[4857]<=16'd4850; ROM2[4857]<=16'd0; ROM3[4857]<=16'd23769; ROM4[4857]<=16'd57273;
ROM1[4858]<=16'd4873; ROM2[4858]<=16'd0; ROM3[4858]<=16'd23779; ROM4[4858]<=16'd57285;
ROM1[4859]<=16'd4865; ROM2[4859]<=16'd0; ROM3[4859]<=16'd23790; ROM4[4859]<=16'd57290;
ROM1[4860]<=16'd4841; ROM2[4860]<=16'd0; ROM3[4860]<=16'd23798; ROM4[4860]<=16'd57287;
ROM1[4861]<=16'd4822; ROM2[4861]<=16'd0; ROM3[4861]<=16'd23793; ROM4[4861]<=16'd57274;
ROM1[4862]<=16'd4819; ROM2[4862]<=16'd0; ROM3[4862]<=16'd23806; ROM4[4862]<=16'd57287;
ROM1[4863]<=16'd4817; ROM2[4863]<=16'd0; ROM3[4863]<=16'd23809; ROM4[4863]<=16'd57292;
ROM1[4864]<=16'd4823; ROM2[4864]<=16'd0; ROM3[4864]<=16'd23789; ROM4[4864]<=16'd57278;
ROM1[4865]<=16'd4852; ROM2[4865]<=16'd0; ROM3[4865]<=16'd23777; ROM4[4865]<=16'd57278;
ROM1[4866]<=16'd4865; ROM2[4866]<=16'd0; ROM3[4866]<=16'd23766; ROM4[4866]<=16'd57273;
ROM1[4867]<=16'd4854; ROM2[4867]<=16'd0; ROM3[4867]<=16'd23767; ROM4[4867]<=16'd57274;
ROM1[4868]<=16'd4833; ROM2[4868]<=16'd0; ROM3[4868]<=16'd23772; ROM4[4868]<=16'd57274;
ROM1[4869]<=16'd4820; ROM2[4869]<=16'd0; ROM3[4869]<=16'd23775; ROM4[4869]<=16'd57270;
ROM1[4870]<=16'd4809; ROM2[4870]<=16'd0; ROM3[4870]<=16'd23786; ROM4[4870]<=16'd57270;
ROM1[4871]<=16'd4801; ROM2[4871]<=16'd0; ROM3[4871]<=16'd23793; ROM4[4871]<=16'd57269;
ROM1[4872]<=16'd4812; ROM2[4872]<=16'd0; ROM3[4872]<=16'd23793; ROM4[4872]<=16'd57274;
ROM1[4873]<=16'd4840; ROM2[4873]<=16'd0; ROM3[4873]<=16'd23787; ROM4[4873]<=16'd57276;
ROM1[4874]<=16'd4870; ROM2[4874]<=16'd0; ROM3[4874]<=16'd23781; ROM4[4874]<=16'd57279;
ROM1[4875]<=16'd4873; ROM2[4875]<=16'd0; ROM3[4875]<=16'd23787; ROM4[4875]<=16'd57283;
ROM1[4876]<=16'd4859; ROM2[4876]<=16'd0; ROM3[4876]<=16'd23795; ROM4[4876]<=16'd57284;
ROM1[4877]<=16'd4851; ROM2[4877]<=16'd0; ROM3[4877]<=16'd23809; ROM4[4877]<=16'd57292;
ROM1[4878]<=16'd4844; ROM2[4878]<=16'd0; ROM3[4878]<=16'd23823; ROM4[4878]<=16'd57300;
ROM1[4879]<=16'd4836; ROM2[4879]<=16'd0; ROM3[4879]<=16'd23834; ROM4[4879]<=16'd57307;
ROM1[4880]<=16'd4834; ROM2[4880]<=16'd0; ROM3[4880]<=16'd23828; ROM4[4880]<=16'd57305;
ROM1[4881]<=16'd4849; ROM2[4881]<=16'd0; ROM3[4881]<=16'd23810; ROM4[4881]<=16'd57297;
ROM1[4882]<=16'd4873; ROM2[4882]<=16'd0; ROM3[4882]<=16'd23787; ROM4[4882]<=16'd57286;
ROM1[4883]<=16'd4865; ROM2[4883]<=16'd0; ROM3[4883]<=16'd23774; ROM4[4883]<=16'd57275;
ROM1[4884]<=16'd4854; ROM2[4884]<=16'd0; ROM3[4884]<=16'd23785; ROM4[4884]<=16'd57279;
ROM1[4885]<=16'd4843; ROM2[4885]<=16'd0; ROM3[4885]<=16'd23799; ROM4[4885]<=16'd57285;
ROM1[4886]<=16'd4822; ROM2[4886]<=16'd0; ROM3[4886]<=16'd23798; ROM4[4886]<=16'd57279;
ROM1[4887]<=16'd4798; ROM2[4887]<=16'd0; ROM3[4887]<=16'd23797; ROM4[4887]<=16'd57273;
ROM1[4888]<=16'd4791; ROM2[4888]<=16'd0; ROM3[4888]<=16'd23794; ROM4[4888]<=16'd57268;
ROM1[4889]<=16'd4808; ROM2[4889]<=16'd0; ROM3[4889]<=16'd23789; ROM4[4889]<=16'd57267;
ROM1[4890]<=16'd4846; ROM2[4890]<=16'd0; ROM3[4890]<=16'd23787; ROM4[4890]<=16'd57275;
ROM1[4891]<=16'd4867; ROM2[4891]<=16'd0; ROM3[4891]<=16'd23784; ROM4[4891]<=16'd57284;
ROM1[4892]<=16'd4870; ROM2[4892]<=16'd0; ROM3[4892]<=16'd23801; ROM4[4892]<=16'd57299;
ROM1[4893]<=16'd4869; ROM2[4893]<=16'd0; ROM3[4893]<=16'd23826; ROM4[4893]<=16'd57315;
ROM1[4894]<=16'd4839; ROM2[4894]<=16'd0; ROM3[4894]<=16'd23822; ROM4[4894]<=16'd57302;
ROM1[4895]<=16'd4814; ROM2[4895]<=16'd0; ROM3[4895]<=16'd23817; ROM4[4895]<=16'd57287;
ROM1[4896]<=16'd4802; ROM2[4896]<=16'd0; ROM3[4896]<=16'd23812; ROM4[4896]<=16'd57279;
ROM1[4897]<=16'd4798; ROM2[4897]<=16'd0; ROM3[4897]<=16'd23800; ROM4[4897]<=16'd57269;
ROM1[4898]<=16'd4845; ROM2[4898]<=16'd0; ROM3[4898]<=16'd23810; ROM4[4898]<=16'd57287;
ROM1[4899]<=16'd4868; ROM2[4899]<=16'd0; ROM3[4899]<=16'd23795; ROM4[4899]<=16'd57283;
ROM1[4900]<=16'd4838; ROM2[4900]<=16'd0; ROM3[4900]<=16'd23779; ROM4[4900]<=16'd57263;
ROM1[4901]<=16'd4817; ROM2[4901]<=16'd0; ROM3[4901]<=16'd23787; ROM4[4901]<=16'd57267;
ROM1[4902]<=16'd4804; ROM2[4902]<=16'd0; ROM3[4902]<=16'd23796; ROM4[4902]<=16'd57270;
ROM1[4903]<=16'd4808; ROM2[4903]<=16'd0; ROM3[4903]<=16'd23817; ROM4[4903]<=16'd57284;
ROM1[4904]<=16'd4812; ROM2[4904]<=16'd0; ROM3[4904]<=16'd23831; ROM4[4904]<=16'd57299;
ROM1[4905]<=16'd4813; ROM2[4905]<=16'd0; ROM3[4905]<=16'd23826; ROM4[4905]<=16'd57291;
ROM1[4906]<=16'd4833; ROM2[4906]<=16'd0; ROM3[4906]<=16'd23812; ROM4[4906]<=16'd57284;
ROM1[4907]<=16'd4869; ROM2[4907]<=16'd0; ROM3[4907]<=16'd23798; ROM4[4907]<=16'd57286;
ROM1[4908]<=16'd4874; ROM2[4908]<=16'd0; ROM3[4908]<=16'd23793; ROM4[4908]<=16'd57284;
ROM1[4909]<=16'd4855; ROM2[4909]<=16'd0; ROM3[4909]<=16'd23798; ROM4[4909]<=16'd57284;
ROM1[4910]<=16'd4839; ROM2[4910]<=16'd0; ROM3[4910]<=16'd23809; ROM4[4910]<=16'd57293;
ROM1[4911]<=16'd4832; ROM2[4911]<=16'd0; ROM3[4911]<=16'd23823; ROM4[4911]<=16'd57301;
ROM1[4912]<=16'd4821; ROM2[4912]<=16'd0; ROM3[4912]<=16'd23833; ROM4[4912]<=16'd57303;
ROM1[4913]<=16'd4812; ROM2[4913]<=16'd0; ROM3[4913]<=16'd23830; ROM4[4913]<=16'd57301;
ROM1[4914]<=16'd4822; ROM2[4914]<=16'd0; ROM3[4914]<=16'd23820; ROM4[4914]<=16'd57293;
ROM1[4915]<=16'd4860; ROM2[4915]<=16'd0; ROM3[4915]<=16'd23814; ROM4[4915]<=16'd57298;
ROM1[4916]<=16'd4894; ROM2[4916]<=16'd0; ROM3[4916]<=16'd23818; ROM4[4916]<=16'd57311;
ROM1[4917]<=16'd4884; ROM2[4917]<=16'd0; ROM3[4917]<=16'd23818; ROM4[4917]<=16'd57308;
ROM1[4918]<=16'd4850; ROM2[4918]<=16'd0; ROM3[4918]<=16'd23811; ROM4[4918]<=16'd57295;
ROM1[4919]<=16'd4830; ROM2[4919]<=16'd0; ROM3[4919]<=16'd23814; ROM4[4919]<=16'd57291;
ROM1[4920]<=16'd4813; ROM2[4920]<=16'd0; ROM3[4920]<=16'd23818; ROM4[4920]<=16'd57290;
ROM1[4921]<=16'd4812; ROM2[4921]<=16'd0; ROM3[4921]<=16'd23826; ROM4[4921]<=16'd57294;
ROM1[4922]<=16'd4824; ROM2[4922]<=16'd0; ROM3[4922]<=16'd23817; ROM4[4922]<=16'd57293;
ROM1[4923]<=16'd4844; ROM2[4923]<=16'd0; ROM3[4923]<=16'd23797; ROM4[4923]<=16'd57283;
ROM1[4924]<=16'd4871; ROM2[4924]<=16'd0; ROM3[4924]<=16'd23786; ROM4[4924]<=16'd57282;
ROM1[4925]<=16'd4874; ROM2[4925]<=16'd0; ROM3[4925]<=16'd23793; ROM4[4925]<=16'd57295;
ROM1[4926]<=16'd4875; ROM2[4926]<=16'd0; ROM3[4926]<=16'd23823; ROM4[4926]<=16'd57314;
ROM1[4927]<=16'd4851; ROM2[4927]<=16'd0; ROM3[4927]<=16'd23828; ROM4[4927]<=16'd57309;
ROM1[4928]<=16'd4814; ROM2[4928]<=16'd0; ROM3[4928]<=16'd23815; ROM4[4928]<=16'd57292;
ROM1[4929]<=16'd4804; ROM2[4929]<=16'd0; ROM3[4929]<=16'd23817; ROM4[4929]<=16'd57288;
ROM1[4930]<=16'd4809; ROM2[4930]<=16'd0; ROM3[4930]<=16'd23808; ROM4[4930]<=16'd57284;
ROM1[4931]<=16'd4837; ROM2[4931]<=16'd0; ROM3[4931]<=16'd23795; ROM4[4931]<=16'd57284;
ROM1[4932]<=16'd4876; ROM2[4932]<=16'd0; ROM3[4932]<=16'd23787; ROM4[4932]<=16'd57286;
ROM1[4933]<=16'd4886; ROM2[4933]<=16'd0; ROM3[4933]<=16'd23785; ROM4[4933]<=16'd57287;
ROM1[4934]<=16'd4862; ROM2[4934]<=16'd0; ROM3[4934]<=16'd23778; ROM4[4934]<=16'd57280;
ROM1[4935]<=16'd4842; ROM2[4935]<=16'd0; ROM3[4935]<=16'd23788; ROM4[4935]<=16'd57277;
ROM1[4936]<=16'd4846; ROM2[4936]<=16'd0; ROM3[4936]<=16'd23812; ROM4[4936]<=16'd57296;
ROM1[4937]<=16'd4823; ROM2[4937]<=16'd0; ROM3[4937]<=16'd23810; ROM4[4937]<=16'd57289;
ROM1[4938]<=16'd4808; ROM2[4938]<=16'd0; ROM3[4938]<=16'd23795; ROM4[4938]<=16'd57271;
ROM1[4939]<=16'd4830; ROM2[4939]<=16'd0; ROM3[4939]<=16'd23789; ROM4[4939]<=16'd57275;
ROM1[4940]<=16'd4859; ROM2[4940]<=16'd0; ROM3[4940]<=16'd23772; ROM4[4940]<=16'd57267;
ROM1[4941]<=16'd4879; ROM2[4941]<=16'd0; ROM3[4941]<=16'd23763; ROM4[4941]<=16'd57270;
ROM1[4942]<=16'd4894; ROM2[4942]<=16'd0; ROM3[4942]<=16'd23789; ROM4[4942]<=16'd57292;
ROM1[4943]<=16'd4872; ROM2[4943]<=16'd0; ROM3[4943]<=16'd23797; ROM4[4943]<=16'd57292;
ROM1[4944]<=16'd4850; ROM2[4944]<=16'd0; ROM3[4944]<=16'd23796; ROM4[4944]<=16'd57285;
ROM1[4945]<=16'd4833; ROM2[4945]<=16'd0; ROM3[4945]<=16'd23806; ROM4[4945]<=16'd57283;
ROM1[4946]<=16'd4823; ROM2[4946]<=16'd0; ROM3[4946]<=16'd23813; ROM4[4946]<=16'd57289;
ROM1[4947]<=16'd4847; ROM2[4947]<=16'd0; ROM3[4947]<=16'd23820; ROM4[4947]<=16'd57300;
ROM1[4948]<=16'd4873; ROM2[4948]<=16'd0; ROM3[4948]<=16'd23808; ROM4[4948]<=16'd57298;
ROM1[4949]<=16'd4892; ROM2[4949]<=16'd0; ROM3[4949]<=16'd23789; ROM4[4949]<=16'd57292;
ROM1[4950]<=16'd4883; ROM2[4950]<=16'd0; ROM3[4950]<=16'd23788; ROM4[4950]<=16'd57290;
ROM1[4951]<=16'd4856; ROM2[4951]<=16'd0; ROM3[4951]<=16'd23786; ROM4[4951]<=16'd57283;
ROM1[4952]<=16'd4844; ROM2[4952]<=16'd0; ROM3[4952]<=16'd23798; ROM4[4952]<=16'd57285;
ROM1[4953]<=16'd4828; ROM2[4953]<=16'd0; ROM3[4953]<=16'd23804; ROM4[4953]<=16'd57283;
ROM1[4954]<=16'd4818; ROM2[4954]<=16'd0; ROM3[4954]<=16'd23806; ROM4[4954]<=16'd57281;
ROM1[4955]<=16'd4825; ROM2[4955]<=16'd0; ROM3[4955]<=16'd23810; ROM4[4955]<=16'd57283;
ROM1[4956]<=16'd4854; ROM2[4956]<=16'd0; ROM3[4956]<=16'd23809; ROM4[4956]<=16'd57291;
ROM1[4957]<=16'd4883; ROM2[4957]<=16'd0; ROM3[4957]<=16'd23795; ROM4[4957]<=16'd57291;
ROM1[4958]<=16'd4867; ROM2[4958]<=16'd0; ROM3[4958]<=16'd23769; ROM4[4958]<=16'd57271;
ROM1[4959]<=16'd4852; ROM2[4959]<=16'd0; ROM3[4959]<=16'd23772; ROM4[4959]<=16'd57272;
ROM1[4960]<=16'd4835; ROM2[4960]<=16'd0; ROM3[4960]<=16'd23777; ROM4[4960]<=16'd57275;
ROM1[4961]<=16'd4825; ROM2[4961]<=16'd0; ROM3[4961]<=16'd23779; ROM4[4961]<=16'd57276;
ROM1[4962]<=16'd4825; ROM2[4962]<=16'd0; ROM3[4962]<=16'd23797; ROM4[4962]<=16'd57288;
ROM1[4963]<=16'd4821; ROM2[4963]<=16'd0; ROM3[4963]<=16'd23796; ROM4[4963]<=16'd57286;
ROM1[4964]<=16'd4832; ROM2[4964]<=16'd0; ROM3[4964]<=16'd23784; ROM4[4964]<=16'd57282;
ROM1[4965]<=16'd4867; ROM2[4965]<=16'd0; ROM3[4965]<=16'd23774; ROM4[4965]<=16'd57286;
ROM1[4966]<=16'd4884; ROM2[4966]<=16'd0; ROM3[4966]<=16'd23768; ROM4[4966]<=16'd57287;
ROM1[4967]<=16'd4869; ROM2[4967]<=16'd0; ROM3[4967]<=16'd23767; ROM4[4967]<=16'd57282;
ROM1[4968]<=16'd4850; ROM2[4968]<=16'd0; ROM3[4968]<=16'd23773; ROM4[4968]<=16'd57278;
ROM1[4969]<=16'd4834; ROM2[4969]<=16'd0; ROM3[4969]<=16'd23785; ROM4[4969]<=16'd57280;
ROM1[4970]<=16'd4821; ROM2[4970]<=16'd0; ROM3[4970]<=16'd23797; ROM4[4970]<=16'd57282;
ROM1[4971]<=16'd4814; ROM2[4971]<=16'd0; ROM3[4971]<=16'd23802; ROM4[4971]<=16'd57283;
ROM1[4972]<=16'd4820; ROM2[4972]<=16'd0; ROM3[4972]<=16'd23791; ROM4[4972]<=16'd57278;
ROM1[4973]<=16'd4844; ROM2[4973]<=16'd0; ROM3[4973]<=16'd23779; ROM4[4973]<=16'd57274;
ROM1[4974]<=16'd4870; ROM2[4974]<=16'd0; ROM3[4974]<=16'd23773; ROM4[4974]<=16'd57276;
ROM1[4975]<=16'd4873; ROM2[4975]<=16'd0; ROM3[4975]<=16'd23778; ROM4[4975]<=16'd57283;
ROM1[4976]<=16'd4862; ROM2[4976]<=16'd0; ROM3[4976]<=16'd23792; ROM4[4976]<=16'd57290;
ROM1[4977]<=16'd4850; ROM2[4977]<=16'd0; ROM3[4977]<=16'd23801; ROM4[4977]<=16'd57289;
ROM1[4978]<=16'd4829; ROM2[4978]<=16'd0; ROM3[4978]<=16'd23797; ROM4[4978]<=16'd57280;
ROM1[4979]<=16'd4810; ROM2[4979]<=16'd0; ROM3[4979]<=16'd23792; ROM4[4979]<=16'd57272;
ROM1[4980]<=16'd4815; ROM2[4980]<=16'd0; ROM3[4980]<=16'd23795; ROM4[4980]<=16'd57273;
ROM1[4981]<=16'd4841; ROM2[4981]<=16'd0; ROM3[4981]<=16'd23789; ROM4[4981]<=16'd57276;
ROM1[4982]<=16'd4871; ROM2[4982]<=16'd0; ROM3[4982]<=16'd23773; ROM4[4982]<=16'd57274;
ROM1[4983]<=16'd4872; ROM2[4983]<=16'd0; ROM3[4983]<=16'd23763; ROM4[4983]<=16'd57266;
ROM1[4984]<=16'd4858; ROM2[4984]<=16'd0; ROM3[4984]<=16'd23765; ROM4[4984]<=16'd57268;
ROM1[4985]<=16'd4855; ROM2[4985]<=16'd0; ROM3[4985]<=16'd23788; ROM4[4985]<=16'd57285;
ROM1[4986]<=16'd4860; ROM2[4986]<=16'd0; ROM3[4986]<=16'd23813; ROM4[4986]<=16'd57306;
ROM1[4987]<=16'd4855; ROM2[4987]<=16'd0; ROM3[4987]<=16'd23832; ROM4[4987]<=16'd57317;
ROM1[4988]<=16'd4856; ROM2[4988]<=16'd0; ROM3[4988]<=16'd23834; ROM4[4988]<=16'd57314;
ROM1[4989]<=16'd4865; ROM2[4989]<=16'd0; ROM3[4989]<=16'd23816; ROM4[4989]<=16'd57306;
ROM1[4990]<=16'd4870; ROM2[4990]<=16'd0; ROM3[4990]<=16'd23784; ROM4[4990]<=16'd57282;
ROM1[4991]<=16'd4868; ROM2[4991]<=16'd0; ROM3[4991]<=16'd23764; ROM4[4991]<=16'd57265;
ROM1[4992]<=16'd4848; ROM2[4992]<=16'd0; ROM3[4992]<=16'd23760; ROM4[4992]<=16'd57258;
ROM1[4993]<=16'd4826; ROM2[4993]<=16'd0; ROM3[4993]<=16'd23766; ROM4[4993]<=16'd57254;
ROM1[4994]<=16'd4830; ROM2[4994]<=16'd0; ROM3[4994]<=16'd23787; ROM4[4994]<=16'd57269;
ROM1[4995]<=16'd4833; ROM2[4995]<=16'd0; ROM3[4995]<=16'd23804; ROM4[4995]<=16'd57284;
ROM1[4996]<=16'd4841; ROM2[4996]<=16'd0; ROM3[4996]<=16'd23822; ROM4[4996]<=16'd57298;
ROM1[4997]<=16'd4842; ROM2[4997]<=16'd0; ROM3[4997]<=16'd23814; ROM4[4997]<=16'd57290;
ROM1[4998]<=16'd4844; ROM2[4998]<=16'd0; ROM3[4998]<=16'd23782; ROM4[4998]<=16'd57267;
ROM1[4999]<=16'd4867; ROM2[4999]<=16'd0; ROM3[4999]<=16'd23770; ROM4[4999]<=16'd57268;
ROM1[5000]<=16'd4862; ROM2[5000]<=16'd0; ROM3[5000]<=16'd23771; ROM4[5000]<=16'd57269;
ROM1[5001]<=16'd4851; ROM2[5001]<=16'd0; ROM3[5001]<=16'd23786; ROM4[5001]<=16'd57275;
ROM1[5002]<=16'd4857; ROM2[5002]<=16'd0; ROM3[5002]<=16'd23815; ROM4[5002]<=16'd57295;
ROM1[5003]<=16'd4840; ROM2[5003]<=16'd0; ROM3[5003]<=16'd23819; ROM4[5003]<=16'd57297;
ROM1[5004]<=16'd4818; ROM2[5004]<=16'd0; ROM3[5004]<=16'd23817; ROM4[5004]<=16'd57288;
ROM1[5005]<=16'd4821; ROM2[5005]<=16'd0; ROM3[5005]<=16'd23811; ROM4[5005]<=16'd57284;
ROM1[5006]<=16'd4852; ROM2[5006]<=16'd0; ROM3[5006]<=16'd23804; ROM4[5006]<=16'd57286;
ROM1[5007]<=16'd4880; ROM2[5007]<=16'd0; ROM3[5007]<=16'd23787; ROM4[5007]<=16'd57279;
ROM1[5008]<=16'd4875; ROM2[5008]<=16'd0; ROM3[5008]<=16'd23777; ROM4[5008]<=16'd57270;
ROM1[5009]<=16'd4860; ROM2[5009]<=16'd0; ROM3[5009]<=16'd23782; ROM4[5009]<=16'd57273;
ROM1[5010]<=16'd4838; ROM2[5010]<=16'd0; ROM3[5010]<=16'd23789; ROM4[5010]<=16'd57273;
ROM1[5011]<=16'd4828; ROM2[5011]<=16'd0; ROM3[5011]<=16'd23799; ROM4[5011]<=16'd57274;
ROM1[5012]<=16'd4818; ROM2[5012]<=16'd0; ROM3[5012]<=16'd23804; ROM4[5012]<=16'd57278;
ROM1[5013]<=16'd4816; ROM2[5013]<=16'd0; ROM3[5013]<=16'd23801; ROM4[5013]<=16'd57274;
ROM1[5014]<=16'd4839; ROM2[5014]<=16'd0; ROM3[5014]<=16'd23798; ROM4[5014]<=16'd57277;
ROM1[5015]<=16'd4879; ROM2[5015]<=16'd0; ROM3[5015]<=16'd23797; ROM4[5015]<=16'd57288;
ROM1[5016]<=16'd4899; ROM2[5016]<=16'd0; ROM3[5016]<=16'd23795; ROM4[5016]<=16'd57292;
ROM1[5017]<=16'd4887; ROM2[5017]<=16'd0; ROM3[5017]<=16'd23797; ROM4[5017]<=16'd57289;
ROM1[5018]<=16'd4868; ROM2[5018]<=16'd0; ROM3[5018]<=16'd23805; ROM4[5018]<=16'd57287;
ROM1[5019]<=16'd4858; ROM2[5019]<=16'd0; ROM3[5019]<=16'd23817; ROM4[5019]<=16'd57287;
ROM1[5020]<=16'd4861; ROM2[5020]<=16'd0; ROM3[5020]<=16'd23839; ROM4[5020]<=16'd57306;
ROM1[5021]<=16'd4859; ROM2[5021]<=16'd0; ROM3[5021]<=16'd23847; ROM4[5021]<=16'd57313;
ROM1[5022]<=16'd4861; ROM2[5022]<=16'd0; ROM3[5022]<=16'd23831; ROM4[5022]<=16'd57301;
ROM1[5023]<=16'd4884; ROM2[5023]<=16'd0; ROM3[5023]<=16'd23812; ROM4[5023]<=16'd57295;
ROM1[5024]<=16'd4888; ROM2[5024]<=16'd0; ROM3[5024]<=16'd23778; ROM4[5024]<=16'd57274;
ROM1[5025]<=16'd4874; ROM2[5025]<=16'd0; ROM3[5025]<=16'd23769; ROM4[5025]<=16'd57265;
ROM1[5026]<=16'd4861; ROM2[5026]<=16'd0; ROM3[5026]<=16'd23779; ROM4[5026]<=16'd57274;
ROM1[5027]<=16'd4840; ROM2[5027]<=16'd0; ROM3[5027]<=16'd23783; ROM4[5027]<=16'd57272;
ROM1[5028]<=16'd4823; ROM2[5028]<=16'd0; ROM3[5028]<=16'd23787; ROM4[5028]<=16'd57271;
ROM1[5029]<=16'd4809; ROM2[5029]<=16'd0; ROM3[5029]<=16'd23789; ROM4[5029]<=16'd57265;
ROM1[5030]<=16'd4818; ROM2[5030]<=16'd0; ROM3[5030]<=16'd23784; ROM4[5030]<=16'd57264;
ROM1[5031]<=16'd4848; ROM2[5031]<=16'd0; ROM3[5031]<=16'd23774; ROM4[5031]<=16'd57266;
ROM1[5032]<=16'd4881; ROM2[5032]<=16'd0; ROM3[5032]<=16'd23769; ROM4[5032]<=16'd57269;
ROM1[5033]<=16'd4886; ROM2[5033]<=16'd0; ROM3[5033]<=16'd23776; ROM4[5033]<=16'd57281;
ROM1[5034]<=16'd4867; ROM2[5034]<=16'd0; ROM3[5034]<=16'd23784; ROM4[5034]<=16'd57284;
ROM1[5035]<=16'd4848; ROM2[5035]<=16'd0; ROM3[5035]<=16'd23794; ROM4[5035]<=16'd57282;
ROM1[5036]<=16'd4838; ROM2[5036]<=16'd0; ROM3[5036]<=16'd23802; ROM4[5036]<=16'd57285;
ROM1[5037]<=16'd4799; ROM2[5037]<=16'd0; ROM3[5037]<=16'd23780; ROM4[5037]<=16'd57257;
ROM1[5038]<=16'd4788; ROM2[5038]<=16'd0; ROM3[5038]<=16'd23771; ROM4[5038]<=16'd57248;
ROM1[5039]<=16'd4810; ROM2[5039]<=16'd0; ROM3[5039]<=16'd23769; ROM4[5039]<=16'd57255;
ROM1[5040]<=16'd4835; ROM2[5040]<=16'd0; ROM3[5040]<=16'd23748; ROM4[5040]<=16'd57251;
ROM1[5041]<=16'd4854; ROM2[5041]<=16'd0; ROM3[5041]<=16'd23746; ROM4[5041]<=16'd57255;
ROM1[5042]<=16'd4848; ROM2[5042]<=16'd0; ROM3[5042]<=16'd23757; ROM4[5042]<=16'd57259;
ROM1[5043]<=16'd4831; ROM2[5043]<=16'd0; ROM3[5043]<=16'd23768; ROM4[5043]<=16'd57262;
ROM1[5044]<=16'd4817; ROM2[5044]<=16'd0; ROM3[5044]<=16'd23775; ROM4[5044]<=16'd57262;
ROM1[5045]<=16'd4807; ROM2[5045]<=16'd0; ROM3[5045]<=16'd23785; ROM4[5045]<=16'd57266;
ROM1[5046]<=16'd4807; ROM2[5046]<=16'd0; ROM3[5046]<=16'd23794; ROM4[5046]<=16'd57272;
ROM1[5047]<=16'd4827; ROM2[5047]<=16'd0; ROM3[5047]<=16'd23799; ROM4[5047]<=16'd57283;
ROM1[5048]<=16'd4864; ROM2[5048]<=16'd0; ROM3[5048]<=16'd23795; ROM4[5048]<=16'd57288;
ROM1[5049]<=16'd4880; ROM2[5049]<=16'd0; ROM3[5049]<=16'd23774; ROM4[5049]<=16'd57278;
ROM1[5050]<=16'd4864; ROM2[5050]<=16'd0; ROM3[5050]<=16'd23762; ROM4[5050]<=16'd57268;
ROM1[5051]<=16'd4848; ROM2[5051]<=16'd0; ROM3[5051]<=16'd23770; ROM4[5051]<=16'd57272;
ROM1[5052]<=16'd4819; ROM2[5052]<=16'd0; ROM3[5052]<=16'd23766; ROM4[5052]<=16'd57265;
ROM1[5053]<=16'd4811; ROM2[5053]<=16'd0; ROM3[5053]<=16'd23777; ROM4[5053]<=16'd57268;
ROM1[5054]<=16'd4818; ROM2[5054]<=16'd0; ROM3[5054]<=16'd23799; ROM4[5054]<=16'd57287;
ROM1[5055]<=16'd4821; ROM2[5055]<=16'd0; ROM3[5055]<=16'd23796; ROM4[5055]<=16'd57283;
ROM1[5056]<=16'd4832; ROM2[5056]<=16'd0; ROM3[5056]<=16'd23772; ROM4[5056]<=16'd57261;
ROM1[5057]<=16'd4854; ROM2[5057]<=16'd0; ROM3[5057]<=16'd23754; ROM4[5057]<=16'd57258;
ROM1[5058]<=16'd4858; ROM2[5058]<=16'd0; ROM3[5058]<=16'd23754; ROM4[5058]<=16'd57261;
ROM1[5059]<=16'd4845; ROM2[5059]<=16'd0; ROM3[5059]<=16'd23759; ROM4[5059]<=16'd57256;
ROM1[5060]<=16'd4837; ROM2[5060]<=16'd0; ROM3[5060]<=16'd23778; ROM4[5060]<=16'd57271;
ROM1[5061]<=16'd4839; ROM2[5061]<=16'd0; ROM3[5061]<=16'd23801; ROM4[5061]<=16'd57286;
ROM1[5062]<=16'd4824; ROM2[5062]<=16'd0; ROM3[5062]<=16'd23811; ROM4[5062]<=16'd57287;
ROM1[5063]<=16'd4808; ROM2[5063]<=16'd0; ROM3[5063]<=16'd23805; ROM4[5063]<=16'd57279;
ROM1[5064]<=16'd4829; ROM2[5064]<=16'd0; ROM3[5064]<=16'd23802; ROM4[5064]<=16'd57279;
ROM1[5065]<=16'd4867; ROM2[5065]<=16'd0; ROM3[5065]<=16'd23789; ROM4[5065]<=16'd57284;
ROM1[5066]<=16'd4883; ROM2[5066]<=16'd0; ROM3[5066]<=16'd23783; ROM4[5066]<=16'd57285;
ROM1[5067]<=16'd4879; ROM2[5067]<=16'd0; ROM3[5067]<=16'd23797; ROM4[5067]<=16'd57292;
ROM1[5068]<=16'd4861; ROM2[5068]<=16'd0; ROM3[5068]<=16'd23808; ROM4[5068]<=16'd57300;
ROM1[5069]<=16'd4838; ROM2[5069]<=16'd0; ROM3[5069]<=16'd23806; ROM4[5069]<=16'd57290;
ROM1[5070]<=16'd4823; ROM2[5070]<=16'd0; ROM3[5070]<=16'd23807; ROM4[5070]<=16'd57284;
ROM1[5071]<=16'd4815; ROM2[5071]<=16'd0; ROM3[5071]<=16'd23803; ROM4[5071]<=16'd57280;
ROM1[5072]<=16'd4826; ROM2[5072]<=16'd0; ROM3[5072]<=16'd23795; ROM4[5072]<=16'd57275;
ROM1[5073]<=16'd4858; ROM2[5073]<=16'd0; ROM3[5073]<=16'd23786; ROM4[5073]<=16'd57277;
ROM1[5074]<=16'd4876; ROM2[5074]<=16'd0; ROM3[5074]<=16'd23762; ROM4[5074]<=16'd57265;
ROM1[5075]<=16'd4861; ROM2[5075]<=16'd0; ROM3[5075]<=16'd23750; ROM4[5075]<=16'd57256;
ROM1[5076]<=16'd4851; ROM2[5076]<=16'd0; ROM3[5076]<=16'd23763; ROM4[5076]<=16'd57262;
ROM1[5077]<=16'd4847; ROM2[5077]<=16'd0; ROM3[5077]<=16'd23781; ROM4[5077]<=16'd57271;
ROM1[5078]<=16'd4829; ROM2[5078]<=16'd0; ROM3[5078]<=16'd23786; ROM4[5078]<=16'd57270;
ROM1[5079]<=16'd4812; ROM2[5079]<=16'd0; ROM3[5079]<=16'd23787; ROM4[5079]<=16'd57269;
ROM1[5080]<=16'd4817; ROM2[5080]<=16'd0; ROM3[5080]<=16'd23785; ROM4[5080]<=16'd57269;
ROM1[5081]<=16'd4836; ROM2[5081]<=16'd0; ROM3[5081]<=16'd23775; ROM4[5081]<=16'd57267;
ROM1[5082]<=16'd4866; ROM2[5082]<=16'd0; ROM3[5082]<=16'd23762; ROM4[5082]<=16'd57261;
ROM1[5083]<=16'd4873; ROM2[5083]<=16'd0; ROM3[5083]<=16'd23762; ROM4[5083]<=16'd57262;
ROM1[5084]<=16'd4861; ROM2[5084]<=16'd0; ROM3[5084]<=16'd23770; ROM4[5084]<=16'd57268;
ROM1[5085]<=16'd4848; ROM2[5085]<=16'd0; ROM3[5085]<=16'd23776; ROM4[5085]<=16'd57271;
ROM1[5086]<=16'd4839; ROM2[5086]<=16'd0; ROM3[5086]<=16'd23786; ROM4[5086]<=16'd57281;
ROM1[5087]<=16'd4807; ROM2[5087]<=16'd0; ROM3[5087]<=16'd23779; ROM4[5087]<=16'd57264;
ROM1[5088]<=16'd4785; ROM2[5088]<=16'd0; ROM3[5088]<=16'd23768; ROM4[5088]<=16'd57243;
ROM1[5089]<=16'd4804; ROM2[5089]<=16'd0; ROM3[5089]<=16'd23770; ROM4[5089]<=16'd57248;
ROM1[5090]<=16'd4832; ROM2[5090]<=16'd0; ROM3[5090]<=16'd23755; ROM4[5090]<=16'd57244;
ROM1[5091]<=16'd4849; ROM2[5091]<=16'd0; ROM3[5091]<=16'd23748; ROM4[5091]<=16'd57248;
ROM1[5092]<=16'd4850; ROM2[5092]<=16'd0; ROM3[5092]<=16'd23758; ROM4[5092]<=16'd57257;
ROM1[5093]<=16'd4823; ROM2[5093]<=16'd0; ROM3[5093]<=16'd23758; ROM4[5093]<=16'd57246;
ROM1[5094]<=16'd4798; ROM2[5094]<=16'd0; ROM3[5094]<=16'd23760; ROM4[5094]<=16'd57240;
ROM1[5095]<=16'd4787; ROM2[5095]<=16'd0; ROM3[5095]<=16'd23773; ROM4[5095]<=16'd57246;
ROM1[5096]<=16'd4779; ROM2[5096]<=16'd0; ROM3[5096]<=16'd23778; ROM4[5096]<=16'd57249;
ROM1[5097]<=16'd4794; ROM2[5097]<=16'd0; ROM3[5097]<=16'd23780; ROM4[5097]<=16'd57257;
ROM1[5098]<=16'd4836; ROM2[5098]<=16'd0; ROM3[5098]<=16'd23783; ROM4[5098]<=16'd57268;
ROM1[5099]<=16'd4868; ROM2[5099]<=16'd0; ROM3[5099]<=16'd23781; ROM4[5099]<=16'd57277;
ROM1[5100]<=16'd4865; ROM2[5100]<=16'd0; ROM3[5100]<=16'd23778; ROM4[5100]<=16'd57277;
ROM1[5101]<=16'd4857; ROM2[5101]<=16'd0; ROM3[5101]<=16'd23791; ROM4[5101]<=16'd57285;
ROM1[5102]<=16'd4855; ROM2[5102]<=16'd0; ROM3[5102]<=16'd23808; ROM4[5102]<=16'd57294;
ROM1[5103]<=16'd4827; ROM2[5103]<=16'd0; ROM3[5103]<=16'd23796; ROM4[5103]<=16'd57277;
ROM1[5104]<=16'd4806; ROM2[5104]<=16'd0; ROM3[5104]<=16'd23788; ROM4[5104]<=16'd57265;
ROM1[5105]<=16'd4816; ROM2[5105]<=16'd0; ROM3[5105]<=16'd23785; ROM4[5105]<=16'd57267;
ROM1[5106]<=16'd4841; ROM2[5106]<=16'd0; ROM3[5106]<=16'd23774; ROM4[5106]<=16'd57268;
ROM1[5107]<=16'd4885; ROM2[5107]<=16'd0; ROM3[5107]<=16'd23773; ROM4[5107]<=16'd57282;
ROM1[5108]<=16'd4881; ROM2[5108]<=16'd0; ROM3[5108]<=16'd23770; ROM4[5108]<=16'd57274;
ROM1[5109]<=16'd4840; ROM2[5109]<=16'd0; ROM3[5109]<=16'd23760; ROM4[5109]<=16'd57253;
ROM1[5110]<=16'd4816; ROM2[5110]<=16'd0; ROM3[5110]<=16'd23766; ROM4[5110]<=16'd57250;
ROM1[5111]<=16'd4808; ROM2[5111]<=16'd0; ROM3[5111]<=16'd23776; ROM4[5111]<=16'd57254;
ROM1[5112]<=16'd4797; ROM2[5112]<=16'd0; ROM3[5112]<=16'd23785; ROM4[5112]<=16'd57260;
ROM1[5113]<=16'd4805; ROM2[5113]<=16'd0; ROM3[5113]<=16'd23799; ROM4[5113]<=16'd57269;
ROM1[5114]<=16'd4824; ROM2[5114]<=16'd0; ROM3[5114]<=16'd23798; ROM4[5114]<=16'd57274;
ROM1[5115]<=16'd4847; ROM2[5115]<=16'd0; ROM3[5115]<=16'd23778; ROM4[5115]<=16'd57272;
ROM1[5116]<=16'd4858; ROM2[5116]<=16'd0; ROM3[5116]<=16'd23768; ROM4[5116]<=16'd57267;
ROM1[5117]<=16'd4849; ROM2[5117]<=16'd0; ROM3[5117]<=16'd23775; ROM4[5117]<=16'd57270;
ROM1[5118]<=16'd4836; ROM2[5118]<=16'd0; ROM3[5118]<=16'd23793; ROM4[5118]<=16'd57279;
ROM1[5119]<=16'd4826; ROM2[5119]<=16'd0; ROM3[5119]<=16'd23807; ROM4[5119]<=16'd57282;
ROM1[5120]<=16'd4815; ROM2[5120]<=16'd0; ROM3[5120]<=16'd23810; ROM4[5120]<=16'd57285;
ROM1[5121]<=16'd4801; ROM2[5121]<=16'd0; ROM3[5121]<=16'd23799; ROM4[5121]<=16'd57277;
ROM1[5122]<=16'd4804; ROM2[5122]<=16'd0; ROM3[5122]<=16'd23782; ROM4[5122]<=16'd57262;
ROM1[5123]<=16'd4836; ROM2[5123]<=16'd0; ROM3[5123]<=16'd23772; ROM4[5123]<=16'd57263;
ROM1[5124]<=16'd4862; ROM2[5124]<=16'd0; ROM3[5124]<=16'd23767; ROM4[5124]<=16'd57264;
ROM1[5125]<=16'd4854; ROM2[5125]<=16'd0; ROM3[5125]<=16'd23774; ROM4[5125]<=16'd57265;
ROM1[5126]<=16'd4832; ROM2[5126]<=16'd0; ROM3[5126]<=16'd23776; ROM4[5126]<=16'd57261;
ROM1[5127]<=16'd4816; ROM2[5127]<=16'd0; ROM3[5127]<=16'd23786; ROM4[5127]<=16'd57263;
ROM1[5128]<=16'd4810; ROM2[5128]<=16'd0; ROM3[5128]<=16'd23802; ROM4[5128]<=16'd57277;
ROM1[5129]<=16'd4809; ROM2[5129]<=16'd0; ROM3[5129]<=16'd23818; ROM4[5129]<=16'd57288;
ROM1[5130]<=16'd4816; ROM2[5130]<=16'd0; ROM3[5130]<=16'd23823; ROM4[5130]<=16'd57295;
ROM1[5131]<=16'd4833; ROM2[5131]<=16'd0; ROM3[5131]<=16'd23805; ROM4[5131]<=16'd57287;
ROM1[5132]<=16'd4864; ROM2[5132]<=16'd0; ROM3[5132]<=16'd23791; ROM4[5132]<=16'd57281;
ROM1[5133]<=16'd4870; ROM2[5133]<=16'd0; ROM3[5133]<=16'd23787; ROM4[5133]<=16'd57283;
ROM1[5134]<=16'd4857; ROM2[5134]<=16'd0; ROM3[5134]<=16'd23793; ROM4[5134]<=16'd57286;
ROM1[5135]<=16'd4837; ROM2[5135]<=16'd0; ROM3[5135]<=16'd23798; ROM4[5135]<=16'd57282;
ROM1[5136]<=16'd4832; ROM2[5136]<=16'd0; ROM3[5136]<=16'd23810; ROM4[5136]<=16'd57288;
ROM1[5137]<=16'd4818; ROM2[5137]<=16'd0; ROM3[5137]<=16'd23814; ROM4[5137]<=16'd57289;
ROM1[5138]<=16'd4814; ROM2[5138]<=16'd0; ROM3[5138]<=16'd23807; ROM4[5138]<=16'd57283;
ROM1[5139]<=16'd4839; ROM2[5139]<=16'd0; ROM3[5139]<=16'd23811; ROM4[5139]<=16'd57289;
ROM1[5140]<=16'd4892; ROM2[5140]<=16'd0; ROM3[5140]<=16'd23819; ROM4[5140]<=16'd57310;
ROM1[5141]<=16'd4916; ROM2[5141]<=16'd0; ROM3[5141]<=16'd23819; ROM4[5141]<=16'd57317;
ROM1[5142]<=16'd4868; ROM2[5142]<=16'd0; ROM3[5142]<=16'd23790; ROM4[5142]<=16'd57279;
ROM1[5143]<=16'd4839; ROM2[5143]<=16'd0; ROM3[5143]<=16'd23781; ROM4[5143]<=16'd57268;
ROM1[5144]<=16'd4824; ROM2[5144]<=16'd0; ROM3[5144]<=16'd23786; ROM4[5144]<=16'd57266;
ROM1[5145]<=16'd4807; ROM2[5145]<=16'd0; ROM3[5145]<=16'd23785; ROM4[5145]<=16'd57260;
ROM1[5146]<=16'd4824; ROM2[5146]<=16'd0; ROM3[5146]<=16'd23806; ROM4[5146]<=16'd57282;
ROM1[5147]<=16'd4838; ROM2[5147]<=16'd0; ROM3[5147]<=16'd23806; ROM4[5147]<=16'd57286;
ROM1[5148]<=16'd4850; ROM2[5148]<=16'd0; ROM3[5148]<=16'd23774; ROM4[5148]<=16'd57265;
ROM1[5149]<=16'd4871; ROM2[5149]<=16'd0; ROM3[5149]<=16'd23762; ROM4[5149]<=16'd57264;
ROM1[5150]<=16'd4870; ROM2[5150]<=16'd0; ROM3[5150]<=16'd23769; ROM4[5150]<=16'd57270;
ROM1[5151]<=16'd4844; ROM2[5151]<=16'd0; ROM3[5151]<=16'd23769; ROM4[5151]<=16'd57262;
ROM1[5152]<=16'd4838; ROM2[5152]<=16'd0; ROM3[5152]<=16'd23792; ROM4[5152]<=16'd57277;
ROM1[5153]<=16'd4808; ROM2[5153]<=16'd0; ROM3[5153]<=16'd23786; ROM4[5153]<=16'd57267;
ROM1[5154]<=16'd4764; ROM2[5154]<=16'd0; ROM3[5154]<=16'd23754; ROM4[5154]<=16'd57237;
ROM1[5155]<=16'd4765; ROM2[5155]<=16'd0; ROM3[5155]<=16'd23747; ROM4[5155]<=16'd57233;
ROM1[5156]<=16'd4784; ROM2[5156]<=16'd0; ROM3[5156]<=16'd23731; ROM4[5156]<=16'd57225;
ROM1[5157]<=16'd4826; ROM2[5157]<=16'd0; ROM3[5157]<=16'd23720; ROM4[5157]<=16'd57224;
ROM1[5158]<=16'd4857; ROM2[5158]<=16'd0; ROM3[5158]<=16'd23744; ROM4[5158]<=16'd57247;
ROM1[5159]<=16'd4850; ROM2[5159]<=16'd0; ROM3[5159]<=16'd23764; ROM4[5159]<=16'd57261;
ROM1[5160]<=16'd4819; ROM2[5160]<=16'd0; ROM3[5160]<=16'd23768; ROM4[5160]<=16'd57256;
ROM1[5161]<=16'd4799; ROM2[5161]<=16'd0; ROM3[5161]<=16'd23773; ROM4[5161]<=16'd57252;
ROM1[5162]<=16'd4788; ROM2[5162]<=16'd0; ROM3[5162]<=16'd23780; ROM4[5162]<=16'd57253;
ROM1[5163]<=16'd4789; ROM2[5163]<=16'd0; ROM3[5163]<=16'd23779; ROM4[5163]<=16'd57254;
ROM1[5164]<=16'd4810; ROM2[5164]<=16'd0; ROM3[5164]<=16'd23773; ROM4[5164]<=16'd57254;
ROM1[5165]<=16'd4839; ROM2[5165]<=16'd0; ROM3[5165]<=16'd23765; ROM4[5165]<=16'd57256;
ROM1[5166]<=16'd4853; ROM2[5166]<=16'd0; ROM3[5166]<=16'd23768; ROM4[5166]<=16'd57261;
ROM1[5167]<=16'd4848; ROM2[5167]<=16'd0; ROM3[5167]<=16'd23777; ROM4[5167]<=16'd57265;
ROM1[5168]<=16'd4836; ROM2[5168]<=16'd0; ROM3[5168]<=16'd23783; ROM4[5168]<=16'd57264;
ROM1[5169]<=16'd4830; ROM2[5169]<=16'd0; ROM3[5169]<=16'd23793; ROM4[5169]<=16'd57268;
ROM1[5170]<=16'd4824; ROM2[5170]<=16'd0; ROM3[5170]<=16'd23798; ROM4[5170]<=16'd57274;
ROM1[5171]<=16'd4812; ROM2[5171]<=16'd0; ROM3[5171]<=16'd23802; ROM4[5171]<=16'd57270;
ROM1[5172]<=16'd4835; ROM2[5172]<=16'd0; ROM3[5172]<=16'd23813; ROM4[5172]<=16'd57284;
ROM1[5173]<=16'd4866; ROM2[5173]<=16'd0; ROM3[5173]<=16'd23807; ROM4[5173]<=16'd57287;
ROM1[5174]<=16'd4881; ROM2[5174]<=16'd0; ROM3[5174]<=16'd23792; ROM4[5174]<=16'd57277;
ROM1[5175]<=16'd4886; ROM2[5175]<=16'd0; ROM3[5175]<=16'd23798; ROM4[5175]<=16'd57281;
ROM1[5176]<=16'd4863; ROM2[5176]<=16'd0; ROM3[5176]<=16'd23800; ROM4[5176]<=16'd57279;
ROM1[5177]<=16'd4838; ROM2[5177]<=16'd0; ROM3[5177]<=16'd23799; ROM4[5177]<=16'd57269;
ROM1[5178]<=16'd4826; ROM2[5178]<=16'd0; ROM3[5178]<=16'd23807; ROM4[5178]<=16'd57278;
ROM1[5179]<=16'd4814; ROM2[5179]<=16'd0; ROM3[5179]<=16'd23811; ROM4[5179]<=16'd57283;
ROM1[5180]<=16'd4818; ROM2[5180]<=16'd0; ROM3[5180]<=16'd23809; ROM4[5180]<=16'd57281;
ROM1[5181]<=16'd4853; ROM2[5181]<=16'd0; ROM3[5181]<=16'd23806; ROM4[5181]<=16'd57295;
ROM1[5182]<=16'd4889; ROM2[5182]<=16'd0; ROM3[5182]<=16'd23800; ROM4[5182]<=16'd57298;
ROM1[5183]<=16'd4888; ROM2[5183]<=16'd0; ROM3[5183]<=16'd23798; ROM4[5183]<=16'd57296;
ROM1[5184]<=16'd4871; ROM2[5184]<=16'd0; ROM3[5184]<=16'd23801; ROM4[5184]<=16'd57294;
ROM1[5185]<=16'd4867; ROM2[5185]<=16'd0; ROM3[5185]<=16'd23816; ROM4[5185]<=16'd57302;
ROM1[5186]<=16'd4868; ROM2[5186]<=16'd0; ROM3[5186]<=16'd23835; ROM4[5186]<=16'd57312;
ROM1[5187]<=16'd4851; ROM2[5187]<=16'd0; ROM3[5187]<=16'd23843; ROM4[5187]<=16'd57311;
ROM1[5188]<=16'd4833; ROM2[5188]<=16'd0; ROM3[5188]<=16'd23827; ROM4[5188]<=16'd57295;
ROM1[5189]<=16'd4826; ROM2[5189]<=16'd0; ROM3[5189]<=16'd23797; ROM4[5189]<=16'd57271;
ROM1[5190]<=16'd4847; ROM2[5190]<=16'd0; ROM3[5190]<=16'd23772; ROM4[5190]<=16'd57256;
ROM1[5191]<=16'd4865; ROM2[5191]<=16'd0; ROM3[5191]<=16'd23763; ROM4[5191]<=16'd57256;
ROM1[5192]<=16'd4867; ROM2[5192]<=16'd0; ROM3[5192]<=16'd23776; ROM4[5192]<=16'd57267;
ROM1[5193]<=16'd4857; ROM2[5193]<=16'd0; ROM3[5193]<=16'd23798; ROM4[5193]<=16'd57277;
ROM1[5194]<=16'd4841; ROM2[5194]<=16'd0; ROM3[5194]<=16'd23806; ROM4[5194]<=16'd57280;
ROM1[5195]<=16'd4819; ROM2[5195]<=16'd0; ROM3[5195]<=16'd23801; ROM4[5195]<=16'd57270;
ROM1[5196]<=16'd4812; ROM2[5196]<=16'd0; ROM3[5196]<=16'd23800; ROM4[5196]<=16'd57270;
ROM1[5197]<=16'd4829; ROM2[5197]<=16'd0; ROM3[5197]<=16'd23800; ROM4[5197]<=16'd57272;
ROM1[5198]<=16'd4870; ROM2[5198]<=16'd0; ROM3[5198]<=16'd23800; ROM4[5198]<=16'd57285;
ROM1[5199]<=16'd4908; ROM2[5199]<=16'd0; ROM3[5199]<=16'd23798; ROM4[5199]<=16'd57295;
ROM1[5200]<=16'd4865; ROM2[5200]<=16'd0; ROM3[5200]<=16'd23761; ROM4[5200]<=16'd57258;
ROM1[5201]<=16'd4823; ROM2[5201]<=16'd0; ROM3[5201]<=16'd23747; ROM4[5201]<=16'd57243;
ROM1[5202]<=16'd4807; ROM2[5202]<=16'd0; ROM3[5202]<=16'd23752; ROM4[5202]<=16'd57242;
ROM1[5203]<=16'd4788; ROM2[5203]<=16'd0; ROM3[5203]<=16'd23755; ROM4[5203]<=16'd57243;
ROM1[5204]<=16'd4798; ROM2[5204]<=16'd0; ROM3[5204]<=16'd23778; ROM4[5204]<=16'd57265;
ROM1[5205]<=16'd4799; ROM2[5205]<=16'd0; ROM3[5205]<=16'd23769; ROM4[5205]<=16'd57253;
ROM1[5206]<=16'd4800; ROM2[5206]<=16'd0; ROM3[5206]<=16'd23741; ROM4[5206]<=16'd57229;
ROM1[5207]<=16'd4831; ROM2[5207]<=16'd0; ROM3[5207]<=16'd23734; ROM4[5207]<=16'd57233;
ROM1[5208]<=16'd4848; ROM2[5208]<=16'd0; ROM3[5208]<=16'd23749; ROM4[5208]<=16'd57249;
ROM1[5209]<=16'd4838; ROM2[5209]<=16'd0; ROM3[5209]<=16'd23768; ROM4[5209]<=16'd57260;
ROM1[5210]<=16'd4822; ROM2[5210]<=16'd0; ROM3[5210]<=16'd23778; ROM4[5210]<=16'd57266;
ROM1[5211]<=16'd4817; ROM2[5211]<=16'd0; ROM3[5211]<=16'd23786; ROM4[5211]<=16'd57271;
ROM1[5212]<=16'd4812; ROM2[5212]<=16'd0; ROM3[5212]<=16'd23800; ROM4[5212]<=16'd57279;
ROM1[5213]<=16'd4806; ROM2[5213]<=16'd0; ROM3[5213]<=16'd23795; ROM4[5213]<=16'd57272;
ROM1[5214]<=16'd4825; ROM2[5214]<=16'd0; ROM3[5214]<=16'd23790; ROM4[5214]<=16'd57273;
ROM1[5215]<=16'd4848; ROM2[5215]<=16'd0; ROM3[5215]<=16'd23772; ROM4[5215]<=16'd57265;
ROM1[5216]<=16'd4845; ROM2[5216]<=16'd0; ROM3[5216]<=16'd23748; ROM4[5216]<=16'd57247;
ROM1[5217]<=16'd4840; ROM2[5217]<=16'd0; ROM3[5217]<=16'd23753; ROM4[5217]<=16'd57254;
ROM1[5218]<=16'd4825; ROM2[5218]<=16'd0; ROM3[5218]<=16'd23765; ROM4[5218]<=16'd57258;
ROM1[5219]<=16'd4806; ROM2[5219]<=16'd0; ROM3[5219]<=16'd23771; ROM4[5219]<=16'd57257;
ROM1[5220]<=16'd4791; ROM2[5220]<=16'd0; ROM3[5220]<=16'd23783; ROM4[5220]<=16'd57264;
ROM1[5221]<=16'd4787; ROM2[5221]<=16'd0; ROM3[5221]<=16'd23793; ROM4[5221]<=16'd57266;
ROM1[5222]<=16'd4802; ROM2[5222]<=16'd0; ROM3[5222]<=16'd23792; ROM4[5222]<=16'd57267;
ROM1[5223]<=16'd4834; ROM2[5223]<=16'd0; ROM3[5223]<=16'd23783; ROM4[5223]<=16'd57267;
ROM1[5224]<=16'd4865; ROM2[5224]<=16'd0; ROM3[5224]<=16'd23783; ROM4[5224]<=16'd57275;
ROM1[5225]<=16'd4864; ROM2[5225]<=16'd0; ROM3[5225]<=16'd23787; ROM4[5225]<=16'd57282;
ROM1[5226]<=16'd4850; ROM2[5226]<=16'd0; ROM3[5226]<=16'd23798; ROM4[5226]<=16'd57287;
ROM1[5227]<=16'd4829; ROM2[5227]<=16'd0; ROM3[5227]<=16'd23803; ROM4[5227]<=16'd57282;
ROM1[5228]<=16'd4815; ROM2[5228]<=16'd0; ROM3[5228]<=16'd23805; ROM4[5228]<=16'd57282;
ROM1[5229]<=16'd4811; ROM2[5229]<=16'd0; ROM3[5229]<=16'd23818; ROM4[5229]<=16'd57291;
ROM1[5230]<=16'd4818; ROM2[5230]<=16'd0; ROM3[5230]<=16'd23817; ROM4[5230]<=16'd57295;
ROM1[5231]<=16'd4844; ROM2[5231]<=16'd0; ROM3[5231]<=16'd23815; ROM4[5231]<=16'd57296;
ROM1[5232]<=16'd4861; ROM2[5232]<=16'd0; ROM3[5232]<=16'd23796; ROM4[5232]<=16'd57282;
ROM1[5233]<=16'd4858; ROM2[5233]<=16'd0; ROM3[5233]<=16'd23791; ROM4[5233]<=16'd57279;
ROM1[5234]<=16'd4829; ROM2[5234]<=16'd0; ROM3[5234]<=16'd23787; ROM4[5234]<=16'd57271;
ROM1[5235]<=16'd4800; ROM2[5235]<=16'd0; ROM3[5235]<=16'd23779; ROM4[5235]<=16'd57261;
ROM1[5236]<=16'd4798; ROM2[5236]<=16'd0; ROM3[5236]<=16'd23786; ROM4[5236]<=16'd57264;
ROM1[5237]<=16'd4783; ROM2[5237]<=16'd0; ROM3[5237]<=16'd23786; ROM4[5237]<=16'd57259;
ROM1[5238]<=16'd4774; ROM2[5238]<=16'd0; ROM3[5238]<=16'd23779; ROM4[5238]<=16'd57253;
ROM1[5239]<=16'd4802; ROM2[5239]<=16'd0; ROM3[5239]<=16'd23785; ROM4[5239]<=16'd57268;
ROM1[5240]<=16'd4838; ROM2[5240]<=16'd0; ROM3[5240]<=16'd23783; ROM4[5240]<=16'd57273;
ROM1[5241]<=16'd4846; ROM2[5241]<=16'd0; ROM3[5241]<=16'd23770; ROM4[5241]<=16'd57265;
ROM1[5242]<=16'd4833; ROM2[5242]<=16'd0; ROM3[5242]<=16'd23767; ROM4[5242]<=16'd57261;
ROM1[5243]<=16'd4813; ROM2[5243]<=16'd0; ROM3[5243]<=16'd23769; ROM4[5243]<=16'd57253;
ROM1[5244]<=16'd4785; ROM2[5244]<=16'd0; ROM3[5244]<=16'd23769; ROM4[5244]<=16'd57247;
ROM1[5245]<=16'd4772; ROM2[5245]<=16'd0; ROM3[5245]<=16'd23775; ROM4[5245]<=16'd57251;
ROM1[5246]<=16'd4771; ROM2[5246]<=16'd0; ROM3[5246]<=16'd23783; ROM4[5246]<=16'd57255;
ROM1[5247]<=16'd4780; ROM2[5247]<=16'd0; ROM3[5247]<=16'd23775; ROM4[5247]<=16'd57252;
ROM1[5248]<=16'd4810; ROM2[5248]<=16'd0; ROM3[5248]<=16'd23761; ROM4[5248]<=16'd57253;
ROM1[5249]<=16'd4833; ROM2[5249]<=16'd0; ROM3[5249]<=16'd23759; ROM4[5249]<=16'd57256;
ROM1[5250]<=16'd4836; ROM2[5250]<=16'd0; ROM3[5250]<=16'd23769; ROM4[5250]<=16'd57262;
ROM1[5251]<=16'd4823; ROM2[5251]<=16'd0; ROM3[5251]<=16'd23778; ROM4[5251]<=16'd57263;
ROM1[5252]<=16'd4829; ROM2[5252]<=16'd0; ROM3[5252]<=16'd23804; ROM4[5252]<=16'd57284;
ROM1[5253]<=16'd4831; ROM2[5253]<=16'd0; ROM3[5253]<=16'd23822; ROM4[5253]<=16'd57298;
ROM1[5254]<=16'd4792; ROM2[5254]<=16'd0; ROM3[5254]<=16'd23801; ROM4[5254]<=16'd57271;
ROM1[5255]<=16'd4770; ROM2[5255]<=16'd0; ROM3[5255]<=16'd23778; ROM4[5255]<=16'd57247;
ROM1[5256]<=16'd4781; ROM2[5256]<=16'd0; ROM3[5256]<=16'd23756; ROM4[5256]<=16'd57235;
ROM1[5257]<=16'd4803; ROM2[5257]<=16'd0; ROM3[5257]<=16'd23734; ROM4[5257]<=16'd57226;
ROM1[5258]<=16'd4816; ROM2[5258]<=16'd0; ROM3[5258]<=16'd23738; ROM4[5258]<=16'd57236;
ROM1[5259]<=16'd4816; ROM2[5259]<=16'd0; ROM3[5259]<=16'd23759; ROM4[5259]<=16'd57250;
ROM1[5260]<=16'd4793; ROM2[5260]<=16'd0; ROM3[5260]<=16'd23762; ROM4[5260]<=16'd57241;
ROM1[5261]<=16'd4773; ROM2[5261]<=16'd0; ROM3[5261]<=16'd23753; ROM4[5261]<=16'd57229;
ROM1[5262]<=16'd4766; ROM2[5262]<=16'd0; ROM3[5262]<=16'd23760; ROM4[5262]<=16'd57237;
ROM1[5263]<=16'd4769; ROM2[5263]<=16'd0; ROM3[5263]<=16'd23764; ROM4[5263]<=16'd57239;
ROM1[5264]<=16'd4785; ROM2[5264]<=16'd0; ROM3[5264]<=16'd23755; ROM4[5264]<=16'd57233;
ROM1[5265]<=16'd4813; ROM2[5265]<=16'd0; ROM3[5265]<=16'd23741; ROM4[5265]<=16'd57228;
ROM1[5266]<=16'd4826; ROM2[5266]<=16'd0; ROM3[5266]<=16'd23737; ROM4[5266]<=16'd57229;
ROM1[5267]<=16'd4818; ROM2[5267]<=16'd0; ROM3[5267]<=16'd23742; ROM4[5267]<=16'd57234;
ROM1[5268]<=16'd4807; ROM2[5268]<=16'd0; ROM3[5268]<=16'd23755; ROM4[5268]<=16'd57240;
ROM1[5269]<=16'd4810; ROM2[5269]<=16'd0; ROM3[5269]<=16'd23781; ROM4[5269]<=16'd57254;
ROM1[5270]<=16'd4802; ROM2[5270]<=16'd0; ROM3[5270]<=16'd23798; ROM4[5270]<=16'd57259;
ROM1[5271]<=16'd4791; ROM2[5271]<=16'd0; ROM3[5271]<=16'd23794; ROM4[5271]<=16'd57255;
ROM1[5272]<=16'd4777; ROM2[5272]<=16'd0; ROM3[5272]<=16'd23765; ROM4[5272]<=16'd57230;
ROM1[5273]<=16'd4782; ROM2[5273]<=16'd0; ROM3[5273]<=16'd23731; ROM4[5273]<=16'd57206;
ROM1[5274]<=16'd4807; ROM2[5274]<=16'd0; ROM3[5274]<=16'd23722; ROM4[5274]<=16'd57207;
ROM1[5275]<=16'd4805; ROM2[5275]<=16'd0; ROM3[5275]<=16'd23730; ROM4[5275]<=16'd57213;
ROM1[5276]<=16'd4803; ROM2[5276]<=16'd0; ROM3[5276]<=16'd23744; ROM4[5276]<=16'd57221;
ROM1[5277]<=16'd4790; ROM2[5277]<=16'd0; ROM3[5277]<=16'd23750; ROM4[5277]<=16'd57221;
ROM1[5278]<=16'd4772; ROM2[5278]<=16'd0; ROM3[5278]<=16'd23749; ROM4[5278]<=16'd57217;
ROM1[5279]<=16'd4762; ROM2[5279]<=16'd0; ROM3[5279]<=16'd23755; ROM4[5279]<=16'd57216;
ROM1[5280]<=16'd4765; ROM2[5280]<=16'd0; ROM3[5280]<=16'd23761; ROM4[5280]<=16'd57220;
ROM1[5281]<=16'd4799; ROM2[5281]<=16'd0; ROM3[5281]<=16'd23763; ROM4[5281]<=16'd57230;
ROM1[5282]<=16'd4836; ROM2[5282]<=16'd0; ROM3[5282]<=16'd23755; ROM4[5282]<=16'd57236;
ROM1[5283]<=16'd4835; ROM2[5283]<=16'd0; ROM3[5283]<=16'd23747; ROM4[5283]<=16'd57231;
ROM1[5284]<=16'd4822; ROM2[5284]<=16'd0; ROM3[5284]<=16'd23759; ROM4[5284]<=16'd57239;
ROM1[5285]<=16'd4819; ROM2[5285]<=16'd0; ROM3[5285]<=16'd23787; ROM4[5285]<=16'd57258;
ROM1[5286]<=16'd4803; ROM2[5286]<=16'd0; ROM3[5286]<=16'd23786; ROM4[5286]<=16'd57250;
ROM1[5287]<=16'd4779; ROM2[5287]<=16'd0; ROM3[5287]<=16'd23775; ROM4[5287]<=16'd57236;
ROM1[5288]<=16'd4781; ROM2[5288]<=16'd0; ROM3[5288]<=16'd23774; ROM4[5288]<=16'd57239;
ROM1[5289]<=16'd4787; ROM2[5289]<=16'd0; ROM3[5289]<=16'd23752; ROM4[5289]<=16'd57230;
ROM1[5290]<=16'd4812; ROM2[5290]<=16'd0; ROM3[5290]<=16'd23738; ROM4[5290]<=16'd57224;
ROM1[5291]<=16'd4831; ROM2[5291]<=16'd0; ROM3[5291]<=16'd23740; ROM4[5291]<=16'd57234;
ROM1[5292]<=16'd4824; ROM2[5292]<=16'd0; ROM3[5292]<=16'd23751; ROM4[5292]<=16'd57239;
ROM1[5293]<=16'd4802; ROM2[5293]<=16'd0; ROM3[5293]<=16'd23759; ROM4[5293]<=16'd57238;
ROM1[5294]<=16'd4796; ROM2[5294]<=16'd0; ROM3[5294]<=16'd23775; ROM4[5294]<=16'd57251;
ROM1[5295]<=16'd4797; ROM2[5295]<=16'd0; ROM3[5295]<=16'd23797; ROM4[5295]<=16'd57270;
ROM1[5296]<=16'd4785; ROM2[5296]<=16'd0; ROM3[5296]<=16'd23790; ROM4[5296]<=16'd57263;
ROM1[5297]<=16'd4789; ROM2[5297]<=16'd0; ROM3[5297]<=16'd23777; ROM4[5297]<=16'd57252;
ROM1[5298]<=16'd4825; ROM2[5298]<=16'd0; ROM3[5298]<=16'd23772; ROM4[5298]<=16'd57259;
ROM1[5299]<=16'd4854; ROM2[5299]<=16'd0; ROM3[5299]<=16'd23766; ROM4[5299]<=16'd57263;
ROM1[5300]<=16'd4851; ROM2[5300]<=16'd0; ROM3[5300]<=16'd23770; ROM4[5300]<=16'd57264;
ROM1[5301]<=16'd4834; ROM2[5301]<=16'd0; ROM3[5301]<=16'd23776; ROM4[5301]<=16'd57266;
ROM1[5302]<=16'd4824; ROM2[5302]<=16'd0; ROM3[5302]<=16'd23793; ROM4[5302]<=16'd57271;
ROM1[5303]<=16'd4820; ROM2[5303]<=16'd0; ROM3[5303]<=16'd23807; ROM4[5303]<=16'd57279;
ROM1[5304]<=16'd4815; ROM2[5304]<=16'd0; ROM3[5304]<=16'd23815; ROM4[5304]<=16'd57289;
ROM1[5305]<=16'd4819; ROM2[5305]<=16'd0; ROM3[5305]<=16'd23814; ROM4[5305]<=16'd57288;
ROM1[5306]<=16'd4829; ROM2[5306]<=16'd0; ROM3[5306]<=16'd23796; ROM4[5306]<=16'd57278;
ROM1[5307]<=16'd4850; ROM2[5307]<=16'd0; ROM3[5307]<=16'd23779; ROM4[5307]<=16'd57271;
ROM1[5308]<=16'd4853; ROM2[5308]<=16'd0; ROM3[5308]<=16'd23771; ROM4[5308]<=16'd57265;
ROM1[5309]<=16'd4841; ROM2[5309]<=16'd0; ROM3[5309]<=16'd23777; ROM4[5309]<=16'd57267;
ROM1[5310]<=16'd4829; ROM2[5310]<=16'd0; ROM3[5310]<=16'd23792; ROM4[5310]<=16'd57272;
ROM1[5311]<=16'd4821; ROM2[5311]<=16'd0; ROM3[5311]<=16'd23798; ROM4[5311]<=16'd57272;
ROM1[5312]<=16'd4809; ROM2[5312]<=16'd0; ROM3[5312]<=16'd23812; ROM4[5312]<=16'd57279;
ROM1[5313]<=16'd4803; ROM2[5313]<=16'd0; ROM3[5313]<=16'd23810; ROM4[5313]<=16'd57276;
ROM1[5314]<=16'd4824; ROM2[5314]<=16'd0; ROM3[5314]<=16'd23800; ROM4[5314]<=16'd57274;
ROM1[5315]<=16'd4844; ROM2[5315]<=16'd0; ROM3[5315]<=16'd23781; ROM4[5315]<=16'd57267;
ROM1[5316]<=16'd4850; ROM2[5316]<=16'd0; ROM3[5316]<=16'd23768; ROM4[5316]<=16'd57258;
ROM1[5317]<=16'd4847; ROM2[5317]<=16'd0; ROM3[5317]<=16'd23779; ROM4[5317]<=16'd57263;
ROM1[5318]<=16'd4833; ROM2[5318]<=16'd0; ROM3[5318]<=16'd23791; ROM4[5318]<=16'd57266;
ROM1[5319]<=16'd4829; ROM2[5319]<=16'd0; ROM3[5319]<=16'd23807; ROM4[5319]<=16'd57276;
ROM1[5320]<=16'd4818; ROM2[5320]<=16'd0; ROM3[5320]<=16'd23814; ROM4[5320]<=16'd57278;
ROM1[5321]<=16'd4803; ROM2[5321]<=16'd0; ROM3[5321]<=16'd23807; ROM4[5321]<=16'd57268;
ROM1[5322]<=16'd4823; ROM2[5322]<=16'd0; ROM3[5322]<=16'd23816; ROM4[5322]<=16'd57280;
ROM1[5323]<=16'd4852; ROM2[5323]<=16'd0; ROM3[5323]<=16'd23804; ROM4[5323]<=16'd57277;
ROM1[5324]<=16'd4861; ROM2[5324]<=16'd0; ROM3[5324]<=16'd23775; ROM4[5324]<=16'd57257;
ROM1[5325]<=16'd4862; ROM2[5325]<=16'd0; ROM3[5325]<=16'd23775; ROM4[5325]<=16'd57259;
ROM1[5326]<=16'd4825; ROM2[5326]<=16'd0; ROM3[5326]<=16'd23759; ROM4[5326]<=16'd57239;
ROM1[5327]<=16'd4799; ROM2[5327]<=16'd0; ROM3[5327]<=16'd23758; ROM4[5327]<=16'd57229;
ROM1[5328]<=16'd4799; ROM2[5328]<=16'd0; ROM3[5328]<=16'd23777; ROM4[5328]<=16'd57246;
ROM1[5329]<=16'd4790; ROM2[5329]<=16'd0; ROM3[5329]<=16'd23779; ROM4[5329]<=16'd57247;
ROM1[5330]<=16'd4804; ROM2[5330]<=16'd0; ROM3[5330]<=16'd23780; ROM4[5330]<=16'd57249;
ROM1[5331]<=16'd4834; ROM2[5331]<=16'd0; ROM3[5331]<=16'd23776; ROM4[5331]<=16'd57259;
ROM1[5332]<=16'd4854; ROM2[5332]<=16'd0; ROM3[5332]<=16'd23758; ROM4[5332]<=16'd57251;
ROM1[5333]<=16'd4859; ROM2[5333]<=16'd0; ROM3[5333]<=16'd23758; ROM4[5333]<=16'd57253;
ROM1[5334]<=16'd4846; ROM2[5334]<=16'd0; ROM3[5334]<=16'd23766; ROM4[5334]<=16'd57255;
ROM1[5335]<=16'd4829; ROM2[5335]<=16'd0; ROM3[5335]<=16'd23771; ROM4[5335]<=16'd57252;
ROM1[5336]<=16'd4828; ROM2[5336]<=16'd0; ROM3[5336]<=16'd23788; ROM4[5336]<=16'd57262;
ROM1[5337]<=16'd4814; ROM2[5337]<=16'd0; ROM3[5337]<=16'd23796; ROM4[5337]<=16'd57265;
ROM1[5338]<=16'd4812; ROM2[5338]<=16'd0; ROM3[5338]<=16'd23795; ROM4[5338]<=16'd57269;
ROM1[5339]<=16'd4837; ROM2[5339]<=16'd0; ROM3[5339]<=16'd23796; ROM4[5339]<=16'd57273;
ROM1[5340]<=16'd4865; ROM2[5340]<=16'd0; ROM3[5340]<=16'd23782; ROM4[5340]<=16'd57267;
ROM1[5341]<=16'd4879; ROM2[5341]<=16'd0; ROM3[5341]<=16'd23779; ROM4[5341]<=16'd57273;
ROM1[5342]<=16'd4869; ROM2[5342]<=16'd0; ROM3[5342]<=16'd23785; ROM4[5342]<=16'd57277;
ROM1[5343]<=16'd4843; ROM2[5343]<=16'd0; ROM3[5343]<=16'd23787; ROM4[5343]<=16'd57271;
ROM1[5344]<=16'd4834; ROM2[5344]<=16'd0; ROM3[5344]<=16'd23799; ROM4[5344]<=16'd57276;
ROM1[5345]<=16'd4822; ROM2[5345]<=16'd0; ROM3[5345]<=16'd23806; ROM4[5345]<=16'd57274;
ROM1[5346]<=16'd4814; ROM2[5346]<=16'd0; ROM3[5346]<=16'd23806; ROM4[5346]<=16'd57271;
ROM1[5347]<=16'd4828; ROM2[5347]<=16'd0; ROM3[5347]<=16'd23800; ROM4[5347]<=16'd57274;
ROM1[5348]<=16'd4862; ROM2[5348]<=16'd0; ROM3[5348]<=16'd23792; ROM4[5348]<=16'd57278;
ROM1[5349]<=16'd4887; ROM2[5349]<=16'd0; ROM3[5349]<=16'd23788; ROM4[5349]<=16'd57284;
ROM1[5350]<=16'd4881; ROM2[5350]<=16'd0; ROM3[5350]<=16'd23794; ROM4[5350]<=16'd57283;
ROM1[5351]<=16'd4862; ROM2[5351]<=16'd0; ROM3[5351]<=16'd23798; ROM4[5351]<=16'd57282;
ROM1[5352]<=16'd4838; ROM2[5352]<=16'd0; ROM3[5352]<=16'd23802; ROM4[5352]<=16'd57280;
ROM1[5353]<=16'd4831; ROM2[5353]<=16'd0; ROM3[5353]<=16'd23813; ROM4[5353]<=16'd57287;
ROM1[5354]<=16'd4832; ROM2[5354]<=16'd0; ROM3[5354]<=16'd23819; ROM4[5354]<=16'd57296;
ROM1[5355]<=16'd4838; ROM2[5355]<=16'd0; ROM3[5355]<=16'd23819; ROM4[5355]<=16'd57295;
ROM1[5356]<=16'd4853; ROM2[5356]<=16'd0; ROM3[5356]<=16'd23805; ROM4[5356]<=16'd57289;
ROM1[5357]<=16'd4879; ROM2[5357]<=16'd0; ROM3[5357]<=16'd23786; ROM4[5357]<=16'd57286;
ROM1[5358]<=16'd4881; ROM2[5358]<=16'd0; ROM3[5358]<=16'd23782; ROM4[5358]<=16'd57284;
ROM1[5359]<=16'd4854; ROM2[5359]<=16'd0; ROM3[5359]<=16'd23782; ROM4[5359]<=16'd57279;
ROM1[5360]<=16'd4833; ROM2[5360]<=16'd0; ROM3[5360]<=16'd23784; ROM4[5360]<=16'd57277;
ROM1[5361]<=16'd4819; ROM2[5361]<=16'd0; ROM3[5361]<=16'd23786; ROM4[5361]<=16'd57273;
ROM1[5362]<=16'd4799; ROM2[5362]<=16'd0; ROM3[5362]<=16'd23786; ROM4[5362]<=16'd57266;
ROM1[5363]<=16'd4801; ROM2[5363]<=16'd0; ROM3[5363]<=16'd23787; ROM4[5363]<=16'd57263;
ROM1[5364]<=16'd4826; ROM2[5364]<=16'd0; ROM3[5364]<=16'd23792; ROM4[5364]<=16'd57272;
ROM1[5365]<=16'd4866; ROM2[5365]<=16'd0; ROM3[5365]<=16'd23797; ROM4[5365]<=16'd57289;
ROM1[5366]<=16'd4867; ROM2[5366]<=16'd0; ROM3[5366]<=16'd23774; ROM4[5366]<=16'd57273;
ROM1[5367]<=16'd4842; ROM2[5367]<=16'd0; ROM3[5367]<=16'd23764; ROM4[5367]<=16'd57257;
ROM1[5368]<=16'd4835; ROM2[5368]<=16'd0; ROM3[5368]<=16'd23781; ROM4[5368]<=16'd57268;
ROM1[5369]<=16'd4816; ROM2[5369]<=16'd0; ROM3[5369]<=16'd23783; ROM4[5369]<=16'd57263;
ROM1[5370]<=16'd4804; ROM2[5370]<=16'd0; ROM3[5370]<=16'd23796; ROM4[5370]<=16'd57271;
ROM1[5371]<=16'd4808; ROM2[5371]<=16'd0; ROM3[5371]<=16'd23811; ROM4[5371]<=16'd57282;
ROM1[5372]<=16'd4824; ROM2[5372]<=16'd0; ROM3[5372]<=16'd23809; ROM4[5372]<=16'd57286;
ROM1[5373]<=16'd4851; ROM2[5373]<=16'd0; ROM3[5373]<=16'd23791; ROM4[5373]<=16'd57279;
ROM1[5374]<=16'd4860; ROM2[5374]<=16'd0; ROM3[5374]<=16'd23767; ROM4[5374]<=16'd57263;
ROM1[5375]<=16'd4860; ROM2[5375]<=16'd0; ROM3[5375]<=16'd23770; ROM4[5375]<=16'd57265;
ROM1[5376]<=16'd4844; ROM2[5376]<=16'd0; ROM3[5376]<=16'd23780; ROM4[5376]<=16'd57265;
ROM1[5377]<=16'd4826; ROM2[5377]<=16'd0; ROM3[5377]<=16'd23786; ROM4[5377]<=16'd57267;
ROM1[5378]<=16'd4821; ROM2[5378]<=16'd0; ROM3[5378]<=16'd23798; ROM4[5378]<=16'd57275;
ROM1[5379]<=16'd4801; ROM2[5379]<=16'd0; ROM3[5379]<=16'd23794; ROM4[5379]<=16'd57266;
ROM1[5380]<=16'd4797; ROM2[5380]<=16'd0; ROM3[5380]<=16'd23782; ROM4[5380]<=16'd57254;
ROM1[5381]<=16'd4821; ROM2[5381]<=16'd0; ROM3[5381]<=16'd23772; ROM4[5381]<=16'd57247;
ROM1[5382]<=16'd4860; ROM2[5382]<=16'd0; ROM3[5382]<=16'd23769; ROM4[5382]<=16'd57257;
ROM1[5383]<=16'd4865; ROM2[5383]<=16'd0; ROM3[5383]<=16'd23771; ROM4[5383]<=16'd57263;
ROM1[5384]<=16'd4854; ROM2[5384]<=16'd0; ROM3[5384]<=16'd23783; ROM4[5384]<=16'd57267;
ROM1[5385]<=16'd4833; ROM2[5385]<=16'd0; ROM3[5385]<=16'd23789; ROM4[5385]<=16'd57265;
ROM1[5386]<=16'd4818; ROM2[5386]<=16'd0; ROM3[5386]<=16'd23792; ROM4[5386]<=16'd57261;
ROM1[5387]<=16'd4811; ROM2[5387]<=16'd0; ROM3[5387]<=16'd23799; ROM4[5387]<=16'd57260;
ROM1[5388]<=16'd4806; ROM2[5388]<=16'd0; ROM3[5388]<=16'd23794; ROM4[5388]<=16'd57254;
ROM1[5389]<=16'd4819; ROM2[5389]<=16'd0; ROM3[5389]<=16'd23787; ROM4[5389]<=16'd57252;
ROM1[5390]<=16'd4854; ROM2[5390]<=16'd0; ROM3[5390]<=16'd23782; ROM4[5390]<=16'd57257;
ROM1[5391]<=16'd4877; ROM2[5391]<=16'd0; ROM3[5391]<=16'd23778; ROM4[5391]<=16'd57261;
ROM1[5392]<=16'd4855; ROM2[5392]<=16'd0; ROM3[5392]<=16'd23768; ROM4[5392]<=16'd57249;
ROM1[5393]<=16'd4841; ROM2[5393]<=16'd0; ROM3[5393]<=16'd23781; ROM4[5393]<=16'd57254;
ROM1[5394]<=16'd4831; ROM2[5394]<=16'd0; ROM3[5394]<=16'd23791; ROM4[5394]<=16'd57260;
ROM1[5395]<=16'd4814; ROM2[5395]<=16'd0; ROM3[5395]<=16'd23801; ROM4[5395]<=16'd57264;
ROM1[5396]<=16'd4820; ROM2[5396]<=16'd0; ROM3[5396]<=16'd23812; ROM4[5396]<=16'd57273;
ROM1[5397]<=16'd4834; ROM2[5397]<=16'd0; ROM3[5397]<=16'd23807; ROM4[5397]<=16'd57269;
ROM1[5398]<=16'd4856; ROM2[5398]<=16'd0; ROM3[5398]<=16'd23789; ROM4[5398]<=16'd57260;
ROM1[5399]<=16'd4871; ROM2[5399]<=16'd0; ROM3[5399]<=16'd23771; ROM4[5399]<=16'd57253;
ROM1[5400]<=16'd4863; ROM2[5400]<=16'd0; ROM3[5400]<=16'd23773; ROM4[5400]<=16'd57254;
ROM1[5401]<=16'd4854; ROM2[5401]<=16'd0; ROM3[5401]<=16'd23787; ROM4[5401]<=16'd57260;
ROM1[5402]<=16'd4845; ROM2[5402]<=16'd0; ROM3[5402]<=16'd23805; ROM4[5402]<=16'd57269;
ROM1[5403]<=16'd4833; ROM2[5403]<=16'd0; ROM3[5403]<=16'd23817; ROM4[5403]<=16'd57275;
ROM1[5404]<=16'd4823; ROM2[5404]<=16'd0; ROM3[5404]<=16'd23819; ROM4[5404]<=16'd57278;
ROM1[5405]<=16'd4825; ROM2[5405]<=16'd0; ROM3[5405]<=16'd23815; ROM4[5405]<=16'd57275;
ROM1[5406]<=16'd4852; ROM2[5406]<=16'd0; ROM3[5406]<=16'd23800; ROM4[5406]<=16'd57273;
ROM1[5407]<=16'd4874; ROM2[5407]<=16'd0; ROM3[5407]<=16'd23776; ROM4[5407]<=16'd57265;
ROM1[5408]<=16'd4881; ROM2[5408]<=16'd0; ROM3[5408]<=16'd23778; ROM4[5408]<=16'd57266;
ROM1[5409]<=16'd4880; ROM2[5409]<=16'd0; ROM3[5409]<=16'd23797; ROM4[5409]<=16'd57281;
ROM1[5410]<=16'd4873; ROM2[5410]<=16'd0; ROM3[5410]<=16'd23820; ROM4[5410]<=16'd57294;
ROM1[5411]<=16'd4848; ROM2[5411]<=16'd0; ROM3[5411]<=16'd23815; ROM4[5411]<=16'd57282;
ROM1[5412]<=16'd4815; ROM2[5412]<=16'd0; ROM3[5412]<=16'd23802; ROM4[5412]<=16'd57264;
ROM1[5413]<=16'd4810; ROM2[5413]<=16'd0; ROM3[5413]<=16'd23794; ROM4[5413]<=16'd57256;
ROM1[5414]<=16'd4825; ROM2[5414]<=16'd0; ROM3[5414]<=16'd23778; ROM4[5414]<=16'd57251;
ROM1[5415]<=16'd4865; ROM2[5415]<=16'd0; ROM3[5415]<=16'd23776; ROM4[5415]<=16'd57256;
ROM1[5416]<=16'd4881; ROM2[5416]<=16'd0; ROM3[5416]<=16'd23775; ROM4[5416]<=16'd57261;
ROM1[5417]<=16'd4879; ROM2[5417]<=16'd0; ROM3[5417]<=16'd23787; ROM4[5417]<=16'd57274;
ROM1[5418]<=16'd4844; ROM2[5418]<=16'd0; ROM3[5418]<=16'd23778; ROM4[5418]<=16'd57256;
ROM1[5419]<=16'd4814; ROM2[5419]<=16'd0; ROM3[5419]<=16'd23769; ROM4[5419]<=16'd57241;
ROM1[5420]<=16'd4809; ROM2[5420]<=16'd0; ROM3[5420]<=16'd23780; ROM4[5420]<=16'd57252;
ROM1[5421]<=16'd4794; ROM2[5421]<=16'd0; ROM3[5421]<=16'd23771; ROM4[5421]<=16'd57243;
ROM1[5422]<=16'd4804; ROM2[5422]<=16'd0; ROM3[5422]<=16'd23763; ROM4[5422]<=16'd57239;
ROM1[5423]<=16'd4855; ROM2[5423]<=16'd0; ROM3[5423]<=16'd23766; ROM4[5423]<=16'd57259;
ROM1[5424]<=16'd4895; ROM2[5424]<=16'd0; ROM3[5424]<=16'd23771; ROM4[5424]<=16'd57272;
ROM1[5425]<=16'd4897; ROM2[5425]<=16'd0; ROM3[5425]<=16'd23780; ROM4[5425]<=16'd57280;
ROM1[5426]<=16'd4892; ROM2[5426]<=16'd0; ROM3[5426]<=16'd23802; ROM4[5426]<=16'd57298;
ROM1[5427]<=16'd4871; ROM2[5427]<=16'd0; ROM3[5427]<=16'd23816; ROM4[5427]<=16'd57299;
ROM1[5428]<=16'd4853; ROM2[5428]<=16'd0; ROM3[5428]<=16'd23818; ROM4[5428]<=16'd57294;
ROM1[5429]<=16'd4844; ROM2[5429]<=16'd0; ROM3[5429]<=16'd23821; ROM4[5429]<=16'd57294;
ROM1[5430]<=16'd4830; ROM2[5430]<=16'd0; ROM3[5430]<=16'd23802; ROM4[5430]<=16'd57273;
ROM1[5431]<=16'd4859; ROM2[5431]<=16'd0; ROM3[5431]<=16'd23788; ROM4[5431]<=16'd57272;
ROM1[5432]<=16'd4896; ROM2[5432]<=16'd0; ROM3[5432]<=16'd23781; ROM4[5432]<=16'd57276;
ROM1[5433]<=16'd4892; ROM2[5433]<=16'd0; ROM3[5433]<=16'd23776; ROM4[5433]<=16'd57269;
ROM1[5434]<=16'd4882; ROM2[5434]<=16'd0; ROM3[5434]<=16'd23790; ROM4[5434]<=16'd57279;
ROM1[5435]<=16'd4857; ROM2[5435]<=16'd0; ROM3[5435]<=16'd23794; ROM4[5435]<=16'd57276;
ROM1[5436]<=16'd4836; ROM2[5436]<=16'd0; ROM3[5436]<=16'd23792; ROM4[5436]<=16'd57271;
ROM1[5437]<=16'd4816; ROM2[5437]<=16'd0; ROM3[5437]<=16'd23788; ROM4[5437]<=16'd57259;
ROM1[5438]<=16'd4824; ROM2[5438]<=16'd0; ROM3[5438]<=16'd23786; ROM4[5438]<=16'd57257;
ROM1[5439]<=16'd4849; ROM2[5439]<=16'd0; ROM3[5439]<=16'd23784; ROM4[5439]<=16'd57259;
ROM1[5440]<=16'd4876; ROM2[5440]<=16'd0; ROM3[5440]<=16'd23774; ROM4[5440]<=16'd57258;
ROM1[5441]<=16'd4894; ROM2[5441]<=16'd0; ROM3[5441]<=16'd23769; ROM4[5441]<=16'd57263;
ROM1[5442]<=16'd4891; ROM2[5442]<=16'd0; ROM3[5442]<=16'd23773; ROM4[5442]<=16'd57268;
ROM1[5443]<=16'd4867; ROM2[5443]<=16'd0; ROM3[5443]<=16'd23775; ROM4[5443]<=16'd57265;
ROM1[5444]<=16'd4849; ROM2[5444]<=16'd0; ROM3[5444]<=16'd23779; ROM4[5444]<=16'd57258;
ROM1[5445]<=16'd4842; ROM2[5445]<=16'd0; ROM3[5445]<=16'd23791; ROM4[5445]<=16'd57263;
ROM1[5446]<=16'd4845; ROM2[5446]<=16'd0; ROM3[5446]<=16'd23803; ROM4[5446]<=16'd57275;
ROM1[5447]<=16'd4861; ROM2[5447]<=16'd0; ROM3[5447]<=16'd23803; ROM4[5447]<=16'd57277;
ROM1[5448]<=16'd4890; ROM2[5448]<=16'd0; ROM3[5448]<=16'd23791; ROM4[5448]<=16'd57276;
ROM1[5449]<=16'd4908; ROM2[5449]<=16'd0; ROM3[5449]<=16'd23779; ROM4[5449]<=16'd57273;
ROM1[5450]<=16'd4892; ROM2[5450]<=16'd0; ROM3[5450]<=16'd23773; ROM4[5450]<=16'd57263;
ROM1[5451]<=16'd4878; ROM2[5451]<=16'd0; ROM3[5451]<=16'd23778; ROM4[5451]<=16'd57265;
ROM1[5452]<=16'd4863; ROM2[5452]<=16'd0; ROM3[5452]<=16'd23782; ROM4[5452]<=16'd57263;
ROM1[5453]<=16'd4840; ROM2[5453]<=16'd0; ROM3[5453]<=16'd23782; ROM4[5453]<=16'd57256;
ROM1[5454]<=16'd4827; ROM2[5454]<=16'd0; ROM3[5454]<=16'd23786; ROM4[5454]<=16'd57258;
ROM1[5455]<=16'd4836; ROM2[5455]<=16'd0; ROM3[5455]<=16'd23789; ROM4[5455]<=16'd57261;
ROM1[5456]<=16'd4858; ROM2[5456]<=16'd0; ROM3[5456]<=16'd23779; ROM4[5456]<=16'd57251;
ROM1[5457]<=16'd4884; ROM2[5457]<=16'd0; ROM3[5457]<=16'd23762; ROM4[5457]<=16'd57247;
ROM1[5458]<=16'd4907; ROM2[5458]<=16'd0; ROM3[5458]<=16'd23778; ROM4[5458]<=16'd57267;
ROM1[5459]<=16'd4893; ROM2[5459]<=16'd0; ROM3[5459]<=16'd23786; ROM4[5459]<=16'd57268;
ROM1[5460]<=16'd4865; ROM2[5460]<=16'd0; ROM3[5460]<=16'd23783; ROM4[5460]<=16'd57261;
ROM1[5461]<=16'd4869; ROM2[5461]<=16'd0; ROM3[5461]<=16'd23803; ROM4[5461]<=16'd57275;
ROM1[5462]<=16'd4857; ROM2[5462]<=16'd0; ROM3[5462]<=16'd23807; ROM4[5462]<=16'd57273;
ROM1[5463]<=16'd4855; ROM2[5463]<=16'd0; ROM3[5463]<=16'd23801; ROM4[5463]<=16'd57271;
ROM1[5464]<=16'd4878; ROM2[5464]<=16'd0; ROM3[5464]<=16'd23798; ROM4[5464]<=16'd57272;
ROM1[5465]<=16'd4897; ROM2[5465]<=16'd0; ROM3[5465]<=16'd23775; ROM4[5465]<=16'd57262;
ROM1[5466]<=16'd4895; ROM2[5466]<=16'd0; ROM3[5466]<=16'd23756; ROM4[5466]<=16'd57247;
ROM1[5467]<=16'd4880; ROM2[5467]<=16'd0; ROM3[5467]<=16'd23761; ROM4[5467]<=16'd57248;
ROM1[5468]<=16'd4873; ROM2[5468]<=16'd0; ROM3[5468]<=16'd23778; ROM4[5468]<=16'd57263;
ROM1[5469]<=16'd4878; ROM2[5469]<=16'd0; ROM3[5469]<=16'd23799; ROM4[5469]<=16'd57275;
ROM1[5470]<=16'd4888; ROM2[5470]<=16'd0; ROM3[5470]<=16'd23825; ROM4[5470]<=16'd57292;
ROM1[5471]<=16'd4869; ROM2[5471]<=16'd0; ROM3[5471]<=16'd23809; ROM4[5471]<=16'd57273;
ROM1[5472]<=16'd4859; ROM2[5472]<=16'd0; ROM3[5472]<=16'd23789; ROM4[5472]<=16'd57255;
ROM1[5473]<=16'd4889; ROM2[5473]<=16'd0; ROM3[5473]<=16'd23782; ROM4[5473]<=16'd57259;
ROM1[5474]<=16'd4898; ROM2[5474]<=16'd0; ROM3[5474]<=16'd23762; ROM4[5474]<=16'd57246;
ROM1[5475]<=16'd4900; ROM2[5475]<=16'd0; ROM3[5475]<=16'd23774; ROM4[5475]<=16'd57255;
ROM1[5476]<=16'd4891; ROM2[5476]<=16'd0; ROM3[5476]<=16'd23780; ROM4[5476]<=16'd57256;
ROM1[5477]<=16'd4863; ROM2[5477]<=16'd0; ROM3[5477]<=16'd23773; ROM4[5477]<=16'd57242;
ROM1[5478]<=16'd4840; ROM2[5478]<=16'd0; ROM3[5478]<=16'd23772; ROM4[5478]<=16'd57236;
ROM1[5479]<=16'd4829; ROM2[5479]<=16'd0; ROM3[5479]<=16'd23777; ROM4[5479]<=16'd57236;
ROM1[5480]<=16'd4844; ROM2[5480]<=16'd0; ROM3[5480]<=16'd23786; ROM4[5480]<=16'd57244;
ROM1[5481]<=16'd4875; ROM2[5481]<=16'd0; ROM3[5481]<=16'd23782; ROM4[5481]<=16'd57249;
ROM1[5482]<=16'd4909; ROM2[5482]<=16'd0; ROM3[5482]<=16'd23772; ROM4[5482]<=16'd57254;
ROM1[5483]<=16'd4903; ROM2[5483]<=16'd0; ROM3[5483]<=16'd23763; ROM4[5483]<=16'd57251;
ROM1[5484]<=16'd4883; ROM2[5484]<=16'd0; ROM3[5484]<=16'd23768; ROM4[5484]<=16'd57250;
ROM1[5485]<=16'd4864; ROM2[5485]<=16'd0; ROM3[5485]<=16'd23774; ROM4[5485]<=16'd57250;
ROM1[5486]<=16'd4847; ROM2[5486]<=16'd0; ROM3[5486]<=16'd23773; ROM4[5486]<=16'd57244;
ROM1[5487]<=16'd4848; ROM2[5487]<=16'd0; ROM3[5487]<=16'd23787; ROM4[5487]<=16'd57254;
ROM1[5488]<=16'd4862; ROM2[5488]<=16'd0; ROM3[5488]<=16'd23799; ROM4[5488]<=16'd57270;
ROM1[5489]<=16'd4873; ROM2[5489]<=16'd0; ROM3[5489]<=16'd23787; ROM4[5489]<=16'd57264;
ROM1[5490]<=16'd4897; ROM2[5490]<=16'd0; ROM3[5490]<=16'd23768; ROM4[5490]<=16'd57253;
ROM1[5491]<=16'd4908; ROM2[5491]<=16'd0; ROM3[5491]<=16'd23762; ROM4[5491]<=16'd57254;
ROM1[5492]<=16'd4892; ROM2[5492]<=16'd0; ROM3[5492]<=16'd23761; ROM4[5492]<=16'd57250;
ROM1[5493]<=16'd4868; ROM2[5493]<=16'd0; ROM3[5493]<=16'd23763; ROM4[5493]<=16'd57243;
ROM1[5494]<=16'd4860; ROM2[5494]<=16'd0; ROM3[5494]<=16'd23774; ROM4[5494]<=16'd57249;
ROM1[5495]<=16'd4853; ROM2[5495]<=16'd0; ROM3[5495]<=16'd23788; ROM4[5495]<=16'd57257;
ROM1[5496]<=16'd4847; ROM2[5496]<=16'd0; ROM3[5496]<=16'd23786; ROM4[5496]<=16'd57255;
ROM1[5497]<=16'd4859; ROM2[5497]<=16'd0; ROM3[5497]<=16'd23780; ROM4[5497]<=16'd57253;
ROM1[5498]<=16'd4887; ROM2[5498]<=16'd0; ROM3[5498]<=16'd23774; ROM4[5498]<=16'd57255;
ROM1[5499]<=16'd4916; ROM2[5499]<=16'd0; ROM3[5499]<=16'd23769; ROM4[5499]<=16'd57260;
ROM1[5500]<=16'd4912; ROM2[5500]<=16'd0; ROM3[5500]<=16'd23770; ROM4[5500]<=16'd57257;
ROM1[5501]<=16'd4911; ROM2[5501]<=16'd0; ROM3[5501]<=16'd23786; ROM4[5501]<=16'd57269;
ROM1[5502]<=16'd4922; ROM2[5502]<=16'd0; ROM3[5502]<=16'd23817; ROM4[5502]<=16'd57292;
ROM1[5503]<=16'd4896; ROM2[5503]<=16'd0; ROM3[5503]<=16'd23808; ROM4[5503]<=16'd57274;
ROM1[5504]<=16'd4881; ROM2[5504]<=16'd0; ROM3[5504]<=16'd23803; ROM4[5504]<=16'd57267;
ROM1[5505]<=16'd4882; ROM2[5505]<=16'd0; ROM3[5505]<=16'd23795; ROM4[5505]<=16'd57260;
ROM1[5506]<=16'd4885; ROM2[5506]<=16'd0; ROM3[5506]<=16'd23762; ROM4[5506]<=16'd57231;
ROM1[5507]<=16'd4920; ROM2[5507]<=16'd0; ROM3[5507]<=16'd23755; ROM4[5507]<=16'd57237;
ROM1[5508]<=16'd4926; ROM2[5508]<=16'd0; ROM3[5508]<=16'd23764; ROM4[5508]<=16'd57243;
ROM1[5509]<=16'd4905; ROM2[5509]<=16'd0; ROM3[5509]<=16'd23767; ROM4[5509]<=16'd57236;
ROM1[5510]<=16'd4879; ROM2[5510]<=16'd0; ROM3[5510]<=16'd23769; ROM4[5510]<=16'd57231;
ROM1[5511]<=16'd4855; ROM2[5511]<=16'd0; ROM3[5511]<=16'd23768; ROM4[5511]<=16'd57225;
ROM1[5512]<=16'd4839; ROM2[5512]<=16'd0; ROM3[5512]<=16'd23764; ROM4[5512]<=16'd57221;
ROM1[5513]<=16'd4836; ROM2[5513]<=16'd0; ROM3[5513]<=16'd23759; ROM4[5513]<=16'd57217;
ROM1[5514]<=16'd4865; ROM2[5514]<=16'd0; ROM3[5514]<=16'd23762; ROM4[5514]<=16'd57230;
ROM1[5515]<=16'd4932; ROM2[5515]<=16'd0; ROM3[5515]<=16'd23777; ROM4[5515]<=16'd57258;
ROM1[5516]<=16'd4930; ROM2[5516]<=16'd0; ROM3[5516]<=16'd23759; ROM4[5516]<=16'd57247;
ROM1[5517]<=16'd4891; ROM2[5517]<=16'd0; ROM3[5517]<=16'd23743; ROM4[5517]<=16'd57231;
ROM1[5518]<=16'd4885; ROM2[5518]<=16'd0; ROM3[5518]<=16'd23759; ROM4[5518]<=16'd57243;
ROM1[5519]<=16'd4867; ROM2[5519]<=16'd0; ROM3[5519]<=16'd23762; ROM4[5519]<=16'd57240;
ROM1[5520]<=16'd4853; ROM2[5520]<=16'd0; ROM3[5520]<=16'd23763; ROM4[5520]<=16'd57239;
ROM1[5521]<=16'd4847; ROM2[5521]<=16'd0; ROM3[5521]<=16'd23766; ROM4[5521]<=16'd57240;
ROM1[5522]<=16'd4852; ROM2[5522]<=16'd0; ROM3[5522]<=16'd23753; ROM4[5522]<=16'd57230;
ROM1[5523]<=16'd4874; ROM2[5523]<=16'd0; ROM3[5523]<=16'd23734; ROM4[5523]<=16'd57224;
ROM1[5524]<=16'd4914; ROM2[5524]<=16'd0; ROM3[5524]<=16'd23743; ROM4[5524]<=16'd57240;
ROM1[5525]<=16'd4928; ROM2[5525]<=16'd0; ROM3[5525]<=16'd23762; ROM4[5525]<=16'd57256;
ROM1[5526]<=16'd4899; ROM2[5526]<=16'd0; ROM3[5526]<=16'd23762; ROM4[5526]<=16'd57246;
ROM1[5527]<=16'd4878; ROM2[5527]<=16'd0; ROM3[5527]<=16'd23764; ROM4[5527]<=16'd57240;
ROM1[5528]<=16'd4869; ROM2[5528]<=16'd0; ROM3[5528]<=16'd23777; ROM4[5528]<=16'd57248;
ROM1[5529]<=16'd4862; ROM2[5529]<=16'd0; ROM3[5529]<=16'd23792; ROM4[5529]<=16'd57257;
ROM1[5530]<=16'd4878; ROM2[5530]<=16'd0; ROM3[5530]<=16'd23804; ROM4[5530]<=16'd57269;
ROM1[5531]<=16'd4910; ROM2[5531]<=16'd0; ROM3[5531]<=16'd23801; ROM4[5531]<=16'd57274;
ROM1[5532]<=16'd4939; ROM2[5532]<=16'd0; ROM3[5532]<=16'd23792; ROM4[5532]<=16'd57270;
ROM1[5533]<=16'd4947; ROM2[5533]<=16'd0; ROM3[5533]<=16'd23798; ROM4[5533]<=16'd57275;
ROM1[5534]<=16'd4926; ROM2[5534]<=16'd0; ROM3[5534]<=16'd23795; ROM4[5534]<=16'd57265;
ROM1[5535]<=16'd4916; ROM2[5535]<=16'd0; ROM3[5535]<=16'd23806; ROM4[5535]<=16'd57270;
ROM1[5536]<=16'd4917; ROM2[5536]<=16'd0; ROM3[5536]<=16'd23826; ROM4[5536]<=16'd57284;
ROM1[5537]<=16'd4887; ROM2[5537]<=16'd0; ROM3[5537]<=16'd23815; ROM4[5537]<=16'd57265;
ROM1[5538]<=16'd4865; ROM2[5538]<=16'd0; ROM3[5538]<=16'd23791; ROM4[5538]<=16'd57245;
ROM1[5539]<=16'd4875; ROM2[5539]<=16'd0; ROM3[5539]<=16'd23774; ROM4[5539]<=16'd57235;
ROM1[5540]<=16'd4905; ROM2[5540]<=16'd0; ROM3[5540]<=16'd23760; ROM4[5540]<=16'd57234;
ROM1[5541]<=16'd4928; ROM2[5541]<=16'd0; ROM3[5541]<=16'd23762; ROM4[5541]<=16'd57244;
ROM1[5542]<=16'd4924; ROM2[5542]<=16'd0; ROM3[5542]<=16'd23779; ROM4[5542]<=16'd57254;
ROM1[5543]<=16'd4896; ROM2[5543]<=16'd0; ROM3[5543]<=16'd23788; ROM4[5543]<=16'd57252;
ROM1[5544]<=16'd4872; ROM2[5544]<=16'd0; ROM3[5544]<=16'd23788; ROM4[5544]<=16'd57244;
ROM1[5545]<=16'd4854; ROM2[5545]<=16'd0; ROM3[5545]<=16'd23794; ROM4[5545]<=16'd57243;
ROM1[5546]<=16'd4848; ROM2[5546]<=16'd0; ROM3[5546]<=16'd23794; ROM4[5546]<=16'd57239;
ROM1[5547]<=16'd4863; ROM2[5547]<=16'd0; ROM3[5547]<=16'd23794; ROM4[5547]<=16'd57242;
ROM1[5548]<=16'd4897; ROM2[5548]<=16'd0; ROM3[5548]<=16'd23791; ROM4[5548]<=16'd57248;
ROM1[5549]<=16'd4906; ROM2[5549]<=16'd0; ROM3[5549]<=16'd23768; ROM4[5549]<=16'd57238;
ROM1[5550]<=16'd4877; ROM2[5550]<=16'd0; ROM3[5550]<=16'd23754; ROM4[5550]<=16'd57226;
ROM1[5551]<=16'd4853; ROM2[5551]<=16'd0; ROM3[5551]<=16'd23757; ROM4[5551]<=16'd57218;
ROM1[5552]<=16'd4832; ROM2[5552]<=16'd0; ROM3[5552]<=16'd23758; ROM4[5552]<=16'd57215;
ROM1[5553]<=16'd4818; ROM2[5553]<=16'd0; ROM3[5553]<=16'd23765; ROM4[5553]<=16'd57218;
ROM1[5554]<=16'd4821; ROM2[5554]<=16'd0; ROM3[5554]<=16'd23785; ROM4[5554]<=16'd57236;
ROM1[5555]<=16'd4826; ROM2[5555]<=16'd0; ROM3[5555]<=16'd23778; ROM4[5555]<=16'd57237;
ROM1[5556]<=16'd4848; ROM2[5556]<=16'd0; ROM3[5556]<=16'd23762; ROM4[5556]<=16'd57236;
ROM1[5557]<=16'd4898; ROM2[5557]<=16'd0; ROM3[5557]<=16'd23765; ROM4[5557]<=16'd57252;
ROM1[5558]<=16'd4923; ROM2[5558]<=16'd0; ROM3[5558]<=16'd23778; ROM4[5558]<=16'd57264;
ROM1[5559]<=16'd4912; ROM2[5559]<=16'd0; ROM3[5559]<=16'd23787; ROM4[5559]<=16'd57270;
ROM1[5560]<=16'd4899; ROM2[5560]<=16'd0; ROM3[5560]<=16'd23802; ROM4[5560]<=16'd57275;
ROM1[5561]<=16'd4885; ROM2[5561]<=16'd0; ROM3[5561]<=16'd23805; ROM4[5561]<=16'd57268;
ROM1[5562]<=16'd4859; ROM2[5562]<=16'd0; ROM3[5562]<=16'd23789; ROM4[5562]<=16'd57250;
ROM1[5563]<=16'd4861; ROM2[5563]<=16'd0; ROM3[5563]<=16'd23788; ROM4[5563]<=16'd57247;
ROM1[5564]<=16'd4886; ROM2[5564]<=16'd0; ROM3[5564]<=16'd23781; ROM4[5564]<=16'd57248;
ROM1[5565]<=16'd4921; ROM2[5565]<=16'd0; ROM3[5565]<=16'd23771; ROM4[5565]<=16'd57254;
ROM1[5566]<=16'd4941; ROM2[5566]<=16'd0; ROM3[5566]<=16'd23779; ROM4[5566]<=16'd57264;
ROM1[5567]<=16'd4929; ROM2[5567]<=16'd0; ROM3[5567]<=16'd23785; ROM4[5567]<=16'd57263;
ROM1[5568]<=16'd4910; ROM2[5568]<=16'd0; ROM3[5568]<=16'd23791; ROM4[5568]<=16'd57262;
ROM1[5569]<=16'd4910; ROM2[5569]<=16'd0; ROM3[5569]<=16'd23813; ROM4[5569]<=16'd57276;
ROM1[5570]<=16'd4919; ROM2[5570]<=16'd0; ROM3[5570]<=16'd23840; ROM4[5570]<=16'd57299;
ROM1[5571]<=16'd4906; ROM2[5571]<=16'd0; ROM3[5571]<=16'd23832; ROM4[5571]<=16'd57294;
ROM1[5572]<=16'd4908; ROM2[5572]<=16'd0; ROM3[5572]<=16'd23818; ROM4[5572]<=16'd57283;
ROM1[5573]<=16'd4923; ROM2[5573]<=16'd0; ROM3[5573]<=16'd23794; ROM4[5573]<=16'd57268;
ROM1[5574]<=16'd4935; ROM2[5574]<=16'd0; ROM3[5574]<=16'd23777; ROM4[5574]<=16'd57259;
ROM1[5575]<=16'd4930; ROM2[5575]<=16'd0; ROM3[5575]<=16'd23782; ROM4[5575]<=16'd57261;
ROM1[5576]<=16'd4913; ROM2[5576]<=16'd0; ROM3[5576]<=16'd23793; ROM4[5576]<=16'd57264;
ROM1[5577]<=16'd4900; ROM2[5577]<=16'd0; ROM3[5577]<=16'd23804; ROM4[5577]<=16'd57265;
ROM1[5578]<=16'd4881; ROM2[5578]<=16'd0; ROM3[5578]<=16'd23803; ROM4[5578]<=16'd57259;
ROM1[5579]<=16'd4881; ROM2[5579]<=16'd0; ROM3[5579]<=16'd23821; ROM4[5579]<=16'd57269;
ROM1[5580]<=16'd4904; ROM2[5580]<=16'd0; ROM3[5580]<=16'd23837; ROM4[5580]<=16'd57287;
ROM1[5581]<=16'd4907; ROM2[5581]<=16'd0; ROM3[5581]<=16'd23813; ROM4[5581]<=16'd57269;
ROM1[5582]<=16'd4905; ROM2[5582]<=16'd0; ROM3[5582]<=16'd23778; ROM4[5582]<=16'd57242;
ROM1[5583]<=16'd4884; ROM2[5583]<=16'd0; ROM3[5583]<=16'd23763; ROM4[5583]<=16'd57223;
ROM1[5584]<=16'd4853; ROM2[5584]<=16'd0; ROM3[5584]<=16'd23762; ROM4[5584]<=16'd57213;
ROM1[5585]<=16'd4849; ROM2[5585]<=16'd0; ROM3[5585]<=16'd23785; ROM4[5585]<=16'd57228;
ROM1[5586]<=16'd4839; ROM2[5586]<=16'd0; ROM3[5586]<=16'd23793; ROM4[5586]<=16'd57232;
ROM1[5587]<=16'd4811; ROM2[5587]<=16'd0; ROM3[5587]<=16'd23783; ROM4[5587]<=16'd57216;
ROM1[5588]<=16'd4806; ROM2[5588]<=16'd0; ROM3[5588]<=16'd23780; ROM4[5588]<=16'd57211;
ROM1[5589]<=16'd4821; ROM2[5589]<=16'd0; ROM3[5589]<=16'd23767; ROM4[5589]<=16'd57209;
ROM1[5590]<=16'd4849; ROM2[5590]<=16'd0; ROM3[5590]<=16'd23752; ROM4[5590]<=16'd57209;
ROM1[5591]<=16'd4869; ROM2[5591]<=16'd0; ROM3[5591]<=16'd23754; ROM4[5591]<=16'd57222;
ROM1[5592]<=16'd4868; ROM2[5592]<=16'd0; ROM3[5592]<=16'd23768; ROM4[5592]<=16'd57233;
ROM1[5593]<=16'd4865; ROM2[5593]<=16'd0; ROM3[5593]<=16'd23793; ROM4[5593]<=16'd57248;
ROM1[5594]<=16'd4839; ROM2[5594]<=16'd0; ROM3[5594]<=16'd23793; ROM4[5594]<=16'd57242;
ROM1[5595]<=16'd4815; ROM2[5595]<=16'd0; ROM3[5595]<=16'd23789; ROM4[5595]<=16'd57234;
ROM1[5596]<=16'd4811; ROM2[5596]<=16'd0; ROM3[5596]<=16'd23781; ROM4[5596]<=16'd57230;
ROM1[5597]<=16'd4822; ROM2[5597]<=16'd0; ROM3[5597]<=16'd23768; ROM4[5597]<=16'd57227;
ROM1[5598]<=16'd4871; ROM2[5598]<=16'd0; ROM3[5598]<=16'd23775; ROM4[5598]<=16'd57245;
ROM1[5599]<=16'd4907; ROM2[5599]<=16'd0; ROM3[5599]<=16'd23778; ROM4[5599]<=16'd57257;
ROM1[5600]<=16'd4904; ROM2[5600]<=16'd0; ROM3[5600]<=16'd23789; ROM4[5600]<=16'd57267;
ROM1[5601]<=16'd4903; ROM2[5601]<=16'd0; ROM3[5601]<=16'd23811; ROM4[5601]<=16'd57284;
ROM1[5602]<=16'd4901; ROM2[5602]<=16'd0; ROM3[5602]<=16'd23822; ROM4[5602]<=16'd57291;
ROM1[5603]<=16'd4879; ROM2[5603]<=16'd0; ROM3[5603]<=16'd23819; ROM4[5603]<=16'd57284;
ROM1[5604]<=16'd4863; ROM2[5604]<=16'd0; ROM3[5604]<=16'd23818; ROM4[5604]<=16'd57281;
ROM1[5605]<=16'd4874; ROM2[5605]<=16'd0; ROM3[5605]<=16'd23817; ROM4[5605]<=16'd57284;
ROM1[5606]<=16'd4893; ROM2[5606]<=16'd0; ROM3[5606]<=16'd23803; ROM4[5606]<=16'd57274;
ROM1[5607]<=16'd4923; ROM2[5607]<=16'd0; ROM3[5607]<=16'd23793; ROM4[5607]<=16'd57279;
ROM1[5608]<=16'd4929; ROM2[5608]<=16'd0; ROM3[5608]<=16'd23795; ROM4[5608]<=16'd57284;
ROM1[5609]<=16'd4897; ROM2[5609]<=16'd0; ROM3[5609]<=16'd23789; ROM4[5609]<=16'd57269;
ROM1[5610]<=16'd4882; ROM2[5610]<=16'd0; ROM3[5610]<=16'd23802; ROM4[5610]<=16'd57277;
ROM1[5611]<=16'd4896; ROM2[5611]<=16'd0; ROM3[5611]<=16'd23834; ROM4[5611]<=16'd57302;
ROM1[5612]<=16'd4878; ROM2[5612]<=16'd0; ROM3[5612]<=16'd23831; ROM4[5612]<=16'd57293;
ROM1[5613]<=16'd4855; ROM2[5613]<=16'd0; ROM3[5613]<=16'd23801; ROM4[5613]<=16'd57264;
ROM1[5614]<=16'd4882; ROM2[5614]<=16'd0; ROM3[5614]<=16'd23796; ROM4[5614]<=16'd57269;
ROM1[5615]<=16'd4919; ROM2[5615]<=16'd0; ROM3[5615]<=16'd23785; ROM4[5615]<=16'd57271;
ROM1[5616]<=16'd4912; ROM2[5616]<=16'd0; ROM3[5616]<=16'd23763; ROM4[5616]<=16'd57252;
ROM1[5617]<=16'd4887; ROM2[5617]<=16'd0; ROM3[5617]<=16'd23763; ROM4[5617]<=16'd57247;
ROM1[5618]<=16'd4856; ROM2[5618]<=16'd0; ROM3[5618]<=16'd23763; ROM4[5618]<=16'd57236;
ROM1[5619]<=16'd4825; ROM2[5619]<=16'd0; ROM3[5619]<=16'd23753; ROM4[5619]<=16'd57218;
ROM1[5620]<=16'd4814; ROM2[5620]<=16'd0; ROM3[5620]<=16'd23756; ROM4[5620]<=16'd57226;
ROM1[5621]<=16'd4824; ROM2[5621]<=16'd0; ROM3[5621]<=16'd23770; ROM4[5621]<=16'd57236;
ROM1[5622]<=16'd4838; ROM2[5622]<=16'd0; ROM3[5622]<=16'd23771; ROM4[5622]<=16'd57239;
ROM1[5623]<=16'd4872; ROM2[5623]<=16'd0; ROM3[5623]<=16'd23759; ROM4[5623]<=16'd57243;
ROM1[5624]<=16'd4897; ROM2[5624]<=16'd0; ROM3[5624]<=16'd23752; ROM4[5624]<=16'd57243;
ROM1[5625]<=16'd4878; ROM2[5625]<=16'd0; ROM3[5625]<=16'd23742; ROM4[5625]<=16'd57234;
ROM1[5626]<=16'd4858; ROM2[5626]<=16'd0; ROM3[5626]<=16'd23745; ROM4[5626]<=16'd57231;
ROM1[5627]<=16'd4846; ROM2[5627]<=16'd0; ROM3[5627]<=16'd23760; ROM4[5627]<=16'd57236;
ROM1[5628]<=16'd4830; ROM2[5628]<=16'd0; ROM3[5628]<=16'd23768; ROM4[5628]<=16'd57243;
ROM1[5629]<=16'd4832; ROM2[5629]<=16'd0; ROM3[5629]<=16'd23786; ROM4[5629]<=16'd57261;
ROM1[5630]<=16'd4849; ROM2[5630]<=16'd0; ROM3[5630]<=16'd23792; ROM4[5630]<=16'd57272;
ROM1[5631]<=16'd4877; ROM2[5631]<=16'd0; ROM3[5631]<=16'd23779; ROM4[5631]<=16'd57273;
ROM1[5632]<=16'd4906; ROM2[5632]<=16'd0; ROM3[5632]<=16'd23771; ROM4[5632]<=16'd57274;
ROM1[5633]<=16'd4916; ROM2[5633]<=16'd0; ROM3[5633]<=16'd23782; ROM4[5633]<=16'd57285;
ROM1[5634]<=16'd4919; ROM2[5634]<=16'd0; ROM3[5634]<=16'd23810; ROM4[5634]<=16'd57308;
ROM1[5635]<=16'd4906; ROM2[5635]<=16'd0; ROM3[5635]<=16'd23826; ROM4[5635]<=16'd57315;
ROM1[5636]<=16'd4881; ROM2[5636]<=16'd0; ROM3[5636]<=16'd23818; ROM4[5636]<=16'd57302;
ROM1[5637]<=16'd4856; ROM2[5637]<=16'd0; ROM3[5637]<=16'd23812; ROM4[5637]<=16'd57290;
ROM1[5638]<=16'd4840; ROM2[5638]<=16'd0; ROM3[5638]<=16'd23798; ROM4[5638]<=16'd57278;
ROM1[5639]<=16'd4847; ROM2[5639]<=16'd0; ROM3[5639]<=16'd23782; ROM4[5639]<=16'd57268;
ROM1[5640]<=16'd4889; ROM2[5640]<=16'd0; ROM3[5640]<=16'd23782; ROM4[5640]<=16'd57272;
ROM1[5641]<=16'd4906; ROM2[5641]<=16'd0; ROM3[5641]<=16'd23785; ROM4[5641]<=16'd57283;
ROM1[5642]<=16'd4873; ROM2[5642]<=16'd0; ROM3[5642]<=16'd23778; ROM4[5642]<=16'd57267;
ROM1[5643]<=16'd4837; ROM2[5643]<=16'd0; ROM3[5643]<=16'd23777; ROM4[5643]<=16'd57251;
ROM1[5644]<=16'd4823; ROM2[5644]<=16'd0; ROM3[5644]<=16'd23783; ROM4[5644]<=16'd57254;
ROM1[5645]<=16'd4813; ROM2[5645]<=16'd0; ROM3[5645]<=16'd23791; ROM4[5645]<=16'd57257;
ROM1[5646]<=16'd4812; ROM2[5646]<=16'd0; ROM3[5646]<=16'd23795; ROM4[5646]<=16'd57259;
ROM1[5647]<=16'd4828; ROM2[5647]<=16'd0; ROM3[5647]<=16'd23796; ROM4[5647]<=16'd57263;
ROM1[5648]<=16'd4852; ROM2[5648]<=16'd0; ROM3[5648]<=16'd23787; ROM4[5648]<=16'd57259;
ROM1[5649]<=16'd4865; ROM2[5649]<=16'd0; ROM3[5649]<=16'd23769; ROM4[5649]<=16'd57250;
ROM1[5650]<=16'd4868; ROM2[5650]<=16'd0; ROM3[5650]<=16'd23779; ROM4[5650]<=16'd57262;
ROM1[5651]<=16'd4864; ROM2[5651]<=16'd0; ROM3[5651]<=16'd23796; ROM4[5651]<=16'd57278;
ROM1[5652]<=16'd4841; ROM2[5652]<=16'd0; ROM3[5652]<=16'd23797; ROM4[5652]<=16'd57274;
ROM1[5653]<=16'd4833; ROM2[5653]<=16'd0; ROM3[5653]<=16'd23810; ROM4[5653]<=16'd57280;
ROM1[5654]<=16'd4832; ROM2[5654]<=16'd0; ROM3[5654]<=16'd23818; ROM4[5654]<=16'd57288;
ROM1[5655]<=16'd4832; ROM2[5655]<=16'd0; ROM3[5655]<=16'd23806; ROM4[5655]<=16'd57277;
ROM1[5656]<=16'd4859; ROM2[5656]<=16'd0; ROM3[5656]<=16'd23793; ROM4[5656]<=16'd57271;
ROM1[5657]<=16'd4890; ROM2[5657]<=16'd0; ROM3[5657]<=16'd23778; ROM4[5657]<=16'd57270;
ROM1[5658]<=16'd4884; ROM2[5658]<=16'd0; ROM3[5658]<=16'd23765; ROM4[5658]<=16'd57260;
ROM1[5659]<=16'd4866; ROM2[5659]<=16'd0; ROM3[5659]<=16'd23770; ROM4[5659]<=16'd57261;
ROM1[5660]<=16'd4853; ROM2[5660]<=16'd0; ROM3[5660]<=16'd23784; ROM4[5660]<=16'd57267;
ROM1[5661]<=16'd4845; ROM2[5661]<=16'd0; ROM3[5661]<=16'd23792; ROM4[5661]<=16'd57271;
ROM1[5662]<=16'd4845; ROM2[5662]<=16'd0; ROM3[5662]<=16'd23809; ROM4[5662]<=16'd57284;
ROM1[5663]<=16'd4847; ROM2[5663]<=16'd0; ROM3[5663]<=16'd23809; ROM4[5663]<=16'd57285;
ROM1[5664]<=16'd4866; ROM2[5664]<=16'd0; ROM3[5664]<=16'd23798; ROM4[5664]<=16'd57288;
ROM1[5665]<=16'd4895; ROM2[5665]<=16'd0; ROM3[5665]<=16'd23784; ROM4[5665]<=16'd57287;
ROM1[5666]<=16'd4890; ROM2[5666]<=16'd0; ROM3[5666]<=16'd23765; ROM4[5666]<=16'd57278;
ROM1[5667]<=16'd4875; ROM2[5667]<=16'd0; ROM3[5667]<=16'd23767; ROM4[5667]<=16'd57279;
ROM1[5668]<=16'd4860; ROM2[5668]<=16'd0; ROM3[5668]<=16'd23780; ROM4[5668]<=16'd57288;
ROM1[5669]<=16'd4846; ROM2[5669]<=16'd0; ROM3[5669]<=16'd23785; ROM4[5669]<=16'd57290;
ROM1[5670]<=16'd4827; ROM2[5670]<=16'd0; ROM3[5670]<=16'd23785; ROM4[5670]<=16'd57282;
ROM1[5671]<=16'd4824; ROM2[5671]<=16'd0; ROM3[5671]<=16'd23789; ROM4[5671]<=16'd57283;
ROM1[5672]<=16'd4853; ROM2[5672]<=16'd0; ROM3[5672]<=16'd23797; ROM4[5672]<=16'd57296;
ROM1[5673]<=16'd4887; ROM2[5673]<=16'd0; ROM3[5673]<=16'd23786; ROM4[5673]<=16'd57293;
ROM1[5674]<=16'd4905; ROM2[5674]<=16'd0; ROM3[5674]<=16'd23771; ROM4[5674]<=16'd57282;
ROM1[5675]<=16'd4899; ROM2[5675]<=16'd0; ROM3[5675]<=16'd23774; ROM4[5675]<=16'd57281;
ROM1[5676]<=16'd4885; ROM2[5676]<=16'd0; ROM3[5676]<=16'd23786; ROM4[5676]<=16'd57284;
ROM1[5677]<=16'd4883; ROM2[5677]<=16'd0; ROM3[5677]<=16'd23812; ROM4[5677]<=16'd57299;
ROM1[5678]<=16'd4866; ROM2[5678]<=16'd0; ROM3[5678]<=16'd23819; ROM4[5678]<=16'd57302;
ROM1[5679]<=16'd4825; ROM2[5679]<=16'd0; ROM3[5679]<=16'd23798; ROM4[5679]<=16'd57275;
ROM1[5680]<=16'd4826; ROM2[5680]<=16'd0; ROM3[5680]<=16'd23785; ROM4[5680]<=16'd57265;
ROM1[5681]<=16'd4858; ROM2[5681]<=16'd0; ROM3[5681]<=16'd23780; ROM4[5681]<=16'd57270;
ROM1[5682]<=16'd4897; ROM2[5682]<=16'd0; ROM3[5682]<=16'd23781; ROM4[5682]<=16'd57278;
ROM1[5683]<=16'd4903; ROM2[5683]<=16'd0; ROM3[5683]<=16'd23784; ROM4[5683]<=16'd57284;
ROM1[5684]<=16'd4870; ROM2[5684]<=16'd0; ROM3[5684]<=16'd23779; ROM4[5684]<=16'd57269;
ROM1[5685]<=16'd4843; ROM2[5685]<=16'd0; ROM3[5685]<=16'd23779; ROM4[5685]<=16'd57261;
ROM1[5686]<=16'd4846; ROM2[5686]<=16'd0; ROM3[5686]<=16'd23796; ROM4[5686]<=16'd57275;
ROM1[5687]<=16'd4840; ROM2[5687]<=16'd0; ROM3[5687]<=16'd23814; ROM4[5687]<=16'd57284;
ROM1[5688]<=16'd4828; ROM2[5688]<=16'd0; ROM3[5688]<=16'd23808; ROM4[5688]<=16'd57275;
ROM1[5689]<=16'd4831; ROM2[5689]<=16'd0; ROM3[5689]<=16'd23788; ROM4[5689]<=16'd57263;
ROM1[5690]<=16'd4838; ROM2[5690]<=16'd0; ROM3[5690]<=16'd23753; ROM4[5690]<=16'd57241;
ROM1[5691]<=16'd4858; ROM2[5691]<=16'd0; ROM3[5691]<=16'd23747; ROM4[5691]<=16'd57246;
ROM1[5692]<=16'd4864; ROM2[5692]<=16'd0; ROM3[5692]<=16'd23766; ROM4[5692]<=16'd57262;
ROM1[5693]<=16'd4844; ROM2[5693]<=16'd0; ROM3[5693]<=16'd23773; ROM4[5693]<=16'd57262;
ROM1[5694]<=16'd4828; ROM2[5694]<=16'd0; ROM3[5694]<=16'd23783; ROM4[5694]<=16'd57266;
ROM1[5695]<=16'd4818; ROM2[5695]<=16'd0; ROM3[5695]<=16'd23795; ROM4[5695]<=16'd57275;
ROM1[5696]<=16'd4822; ROM2[5696]<=16'd0; ROM3[5696]<=16'd23802; ROM4[5696]<=16'd57285;
ROM1[5697]<=16'd4849; ROM2[5697]<=16'd0; ROM3[5697]<=16'd23804; ROM4[5697]<=16'd57291;
ROM1[5698]<=16'd4883; ROM2[5698]<=16'd0; ROM3[5698]<=16'd23796; ROM4[5698]<=16'd57292;
ROM1[5699]<=16'd4900; ROM2[5699]<=16'd0; ROM3[5699]<=16'd23787; ROM4[5699]<=16'd57294;
ROM1[5700]<=16'd4885; ROM2[5700]<=16'd0; ROM3[5700]<=16'd23786; ROM4[5700]<=16'd57292;
ROM1[5701]<=16'd4853; ROM2[5701]<=16'd0; ROM3[5701]<=16'd23784; ROM4[5701]<=16'd57283;
ROM1[5702]<=16'd4844; ROM2[5702]<=16'd0; ROM3[5702]<=16'd23797; ROM4[5702]<=16'd57289;
ROM1[5703]<=16'd4832; ROM2[5703]<=16'd0; ROM3[5703]<=16'd23800; ROM4[5703]<=16'd57282;
ROM1[5704]<=16'd4806; ROM2[5704]<=16'd0; ROM3[5704]<=16'd23789; ROM4[5704]<=16'd57264;
ROM1[5705]<=16'd4807; ROM2[5705]<=16'd0; ROM3[5705]<=16'd23785; ROM4[5705]<=16'd57261;
ROM1[5706]<=16'd4829; ROM2[5706]<=16'd0; ROM3[5706]<=16'd23769; ROM4[5706]<=16'd57256;
ROM1[5707]<=16'd4858; ROM2[5707]<=16'd0; ROM3[5707]<=16'd23757; ROM4[5707]<=16'd57255;
ROM1[5708]<=16'd4856; ROM2[5708]<=16'd0; ROM3[5708]<=16'd23747; ROM4[5708]<=16'd57250;
ROM1[5709]<=16'd4837; ROM2[5709]<=16'd0; ROM3[5709]<=16'd23748; ROM4[5709]<=16'd57250;
ROM1[5710]<=16'd4828; ROM2[5710]<=16'd0; ROM3[5710]<=16'd23768; ROM4[5710]<=16'd57261;
ROM1[5711]<=16'd4815; ROM2[5711]<=16'd0; ROM3[5711]<=16'd23773; ROM4[5711]<=16'd57260;
ROM1[5712]<=16'd4806; ROM2[5712]<=16'd0; ROM3[5712]<=16'd23782; ROM4[5712]<=16'd57265;
ROM1[5713]<=16'd4818; ROM2[5713]<=16'd0; ROM3[5713]<=16'd23793; ROM4[5713]<=16'd57277;
ROM1[5714]<=16'd4835; ROM2[5714]<=16'd0; ROM3[5714]<=16'd23785; ROM4[5714]<=16'd57273;
ROM1[5715]<=16'd4853; ROM2[5715]<=16'd0; ROM3[5715]<=16'd23762; ROM4[5715]<=16'd57263;
ROM1[5716]<=16'd4857; ROM2[5716]<=16'd0; ROM3[5716]<=16'd23750; ROM4[5716]<=16'd57259;
ROM1[5717]<=16'd4838; ROM2[5717]<=16'd0; ROM3[5717]<=16'd23747; ROM4[5717]<=16'd57254;
ROM1[5718]<=16'd4814; ROM2[5718]<=16'd0; ROM3[5718]<=16'd23747; ROM4[5718]<=16'd57249;
ROM1[5719]<=16'd4814; ROM2[5719]<=16'd0; ROM3[5719]<=16'd23759; ROM4[5719]<=16'd57261;
ROM1[5720]<=16'd4812; ROM2[5720]<=16'd0; ROM3[5720]<=16'd23780; ROM4[5720]<=16'd57275;
ROM1[5721]<=16'd4812; ROM2[5721]<=16'd0; ROM3[5721]<=16'd23788; ROM4[5721]<=16'd57279;
ROM1[5722]<=16'd4817; ROM2[5722]<=16'd0; ROM3[5722]<=16'd23775; ROM4[5722]<=16'd57271;
ROM1[5723]<=16'd4838; ROM2[5723]<=16'd0; ROM3[5723]<=16'd23754; ROM4[5723]<=16'd57259;
ROM1[5724]<=16'd4855; ROM2[5724]<=16'd0; ROM3[5724]<=16'd23737; ROM4[5724]<=16'd57253;
ROM1[5725]<=16'd4837; ROM2[5725]<=16'd0; ROM3[5725]<=16'd23727; ROM4[5725]<=16'd57245;
ROM1[5726]<=16'd4823; ROM2[5726]<=16'd0; ROM3[5726]<=16'd23742; ROM4[5726]<=16'd57254;
ROM1[5727]<=16'd4826; ROM2[5727]<=16'd0; ROM3[5727]<=16'd23772; ROM4[5727]<=16'd57272;
ROM1[5728]<=16'd4810; ROM2[5728]<=16'd0; ROM3[5728]<=16'd23781; ROM4[5728]<=16'd57268;
ROM1[5729]<=16'd4800; ROM2[5729]<=16'd0; ROM3[5729]<=16'd23782; ROM4[5729]<=16'd57261;
ROM1[5730]<=16'd4814; ROM2[5730]<=16'd0; ROM3[5730]<=16'd23786; ROM4[5730]<=16'd57268;
ROM1[5731]<=16'd4839; ROM2[5731]<=16'd0; ROM3[5731]<=16'd23784; ROM4[5731]<=16'd57274;
ROM1[5732]<=16'd4857; ROM2[5732]<=16'd0; ROM3[5732]<=16'd23772; ROM4[5732]<=16'd57268;
ROM1[5733]<=16'd4850; ROM2[5733]<=16'd0; ROM3[5733]<=16'd23767; ROM4[5733]<=16'd57265;
ROM1[5734]<=16'd4834; ROM2[5734]<=16'd0; ROM3[5734]<=16'd23771; ROM4[5734]<=16'd57263;
ROM1[5735]<=16'd4826; ROM2[5735]<=16'd0; ROM3[5735]<=16'd23786; ROM4[5735]<=16'd57271;
ROM1[5736]<=16'd4832; ROM2[5736]<=16'd0; ROM3[5736]<=16'd23808; ROM4[5736]<=16'd57290;
ROM1[5737]<=16'd4819; ROM2[5737]<=16'd0; ROM3[5737]<=16'd23815; ROM4[5737]<=16'd57288;
ROM1[5738]<=16'd4807; ROM2[5738]<=16'd0; ROM3[5738]<=16'd23803; ROM4[5738]<=16'd57278;
ROM1[5739]<=16'd4818; ROM2[5739]<=16'd0; ROM3[5739]<=16'd23786; ROM4[5739]<=16'd57269;
ROM1[5740]<=16'd4850; ROM2[5740]<=16'd0; ROM3[5740]<=16'd23773; ROM4[5740]<=16'd57268;
ROM1[5741]<=16'd4865; ROM2[5741]<=16'd0; ROM3[5741]<=16'd23773; ROM4[5741]<=16'd57275;
ROM1[5742]<=16'd4857; ROM2[5742]<=16'd0; ROM3[5742]<=16'd23782; ROM4[5742]<=16'd57280;
ROM1[5743]<=16'd4833; ROM2[5743]<=16'd0; ROM3[5743]<=16'd23781; ROM4[5743]<=16'd57275;
ROM1[5744]<=16'd4813; ROM2[5744]<=16'd0; ROM3[5744]<=16'd23782; ROM4[5744]<=16'd57274;
ROM1[5745]<=16'd4807; ROM2[5745]<=16'd0; ROM3[5745]<=16'd23794; ROM4[5745]<=16'd57283;
ROM1[5746]<=16'd4803; ROM2[5746]<=16'd0; ROM3[5746]<=16'd23795; ROM4[5746]<=16'd57278;
ROM1[5747]<=16'd4822; ROM2[5747]<=16'd0; ROM3[5747]<=16'd23796; ROM4[5747]<=16'd57286;
ROM1[5748]<=16'd4846; ROM2[5748]<=16'd0; ROM3[5748]<=16'd23781; ROM4[5748]<=16'd57279;
ROM1[5749]<=16'd4850; ROM2[5749]<=16'd0; ROM3[5749]<=16'd23755; ROM4[5749]<=16'd57261;
ROM1[5750]<=16'd4852; ROM2[5750]<=16'd0; ROM3[5750]<=16'd23770; ROM4[5750]<=16'd57276;
ROM1[5751]<=16'd4820; ROM2[5751]<=16'd0; ROM3[5751]<=16'd23768; ROM4[5751]<=16'd57267;
ROM1[5752]<=16'd4784; ROM2[5752]<=16'd0; ROM3[5752]<=16'd23757; ROM4[5752]<=16'd57251;
ROM1[5753]<=16'd4777; ROM2[5753]<=16'd0; ROM3[5753]<=16'd23771; ROM4[5753]<=16'd57261;
ROM1[5754]<=16'd4771; ROM2[5754]<=16'd0; ROM3[5754]<=16'd23778; ROM4[5754]<=16'd57265;
ROM1[5755]<=16'd4785; ROM2[5755]<=16'd0; ROM3[5755]<=16'd23783; ROM4[5755]<=16'd57270;
ROM1[5756]<=16'd4815; ROM2[5756]<=16'd0; ROM3[5756]<=16'd23780; ROM4[5756]<=16'd57274;
ROM1[5757]<=16'd4845; ROM2[5757]<=16'd0; ROM3[5757]<=16'd23767; ROM4[5757]<=16'd57277;
ROM1[5758]<=16'd4841; ROM2[5758]<=16'd0; ROM3[5758]<=16'd23759; ROM4[5758]<=16'd57271;
ROM1[5759]<=16'd4827; ROM2[5759]<=16'd0; ROM3[5759]<=16'd23761; ROM4[5759]<=16'd57266;
ROM1[5760]<=16'd4817; ROM2[5760]<=16'd0; ROM3[5760]<=16'd23773; ROM4[5760]<=16'd57278;
ROM1[5761]<=16'd4808; ROM2[5761]<=16'd0; ROM3[5761]<=16'd23783; ROM4[5761]<=16'd57279;
ROM1[5762]<=16'd4793; ROM2[5762]<=16'd0; ROM3[5762]<=16'd23784; ROM4[5762]<=16'd57273;
ROM1[5763]<=16'd4785; ROM2[5763]<=16'd0; ROM3[5763]<=16'd23773; ROM4[5763]<=16'd57265;
ROM1[5764]<=16'd4797; ROM2[5764]<=16'd0; ROM3[5764]<=16'd23760; ROM4[5764]<=16'd57256;
ROM1[5765]<=16'd4828; ROM2[5765]<=16'd0; ROM3[5765]<=16'd23749; ROM4[5765]<=16'd57254;
ROM1[5766]<=16'd4831; ROM2[5766]<=16'd0; ROM3[5766]<=16'd23738; ROM4[5766]<=16'd57251;
ROM1[5767]<=16'd4819; ROM2[5767]<=16'd0; ROM3[5767]<=16'd23744; ROM4[5767]<=16'd57253;
ROM1[5768]<=16'd4809; ROM2[5768]<=16'd0; ROM3[5768]<=16'd23752; ROM4[5768]<=16'd57255;
ROM1[5769]<=16'd4792; ROM2[5769]<=16'd0; ROM3[5769]<=16'd23751; ROM4[5769]<=16'd57248;
ROM1[5770]<=16'd4779; ROM2[5770]<=16'd0; ROM3[5770]<=16'd23759; ROM4[5770]<=16'd57251;
ROM1[5771]<=16'd4777; ROM2[5771]<=16'd0; ROM3[5771]<=16'd23764; ROM4[5771]<=16'd57257;
ROM1[5772]<=16'd4814; ROM2[5772]<=16'd0; ROM3[5772]<=16'd23782; ROM4[5772]<=16'd57280;
ROM1[5773]<=16'd4853; ROM2[5773]<=16'd0; ROM3[5773]<=16'd23776; ROM4[5773]<=16'd57288;
ROM1[5774]<=16'd4853; ROM2[5774]<=16'd0; ROM3[5774]<=16'd23750; ROM4[5774]<=16'd57270;
ROM1[5775]<=16'd4838; ROM2[5775]<=16'd0; ROM3[5775]<=16'd23743; ROM4[5775]<=16'd57262;
ROM1[5776]<=16'd4822; ROM2[5776]<=16'd0; ROM3[5776]<=16'd23750; ROM4[5776]<=16'd57263;
ROM1[5777]<=16'd4799; ROM2[5777]<=16'd0; ROM3[5777]<=16'd23753; ROM4[5777]<=16'd57255;
ROM1[5778]<=16'd4786; ROM2[5778]<=16'd0; ROM3[5778]<=16'd23755; ROM4[5778]<=16'd57253;
ROM1[5779]<=16'd4796; ROM2[5779]<=16'd0; ROM3[5779]<=16'd23774; ROM4[5779]<=16'd57271;
ROM1[5780]<=16'd4794; ROM2[5780]<=16'd0; ROM3[5780]<=16'd23764; ROM4[5780]<=16'd57265;
ROM1[5781]<=16'd4806; ROM2[5781]<=16'd0; ROM3[5781]<=16'd23743; ROM4[5781]<=16'd57253;
ROM1[5782]<=16'd4846; ROM2[5782]<=16'd0; ROM3[5782]<=16'd23745; ROM4[5782]<=16'd57263;
ROM1[5783]<=16'd4849; ROM2[5783]<=16'd0; ROM3[5783]<=16'd23755; ROM4[5783]<=16'd57269;
ROM1[5784]<=16'd4839; ROM2[5784]<=16'd0; ROM3[5784]<=16'd23766; ROM4[5784]<=16'd57275;
ROM1[5785]<=16'd4835; ROM2[5785]<=16'd0; ROM3[5785]<=16'd23785; ROM4[5785]<=16'd57286;
ROM1[5786]<=16'd4823; ROM2[5786]<=16'd0; ROM3[5786]<=16'd23796; ROM4[5786]<=16'd57290;
ROM1[5787]<=16'd4803; ROM2[5787]<=16'd0; ROM3[5787]<=16'd23802; ROM4[5787]<=16'd57286;
ROM1[5788]<=16'd4812; ROM2[5788]<=16'd0; ROM3[5788]<=16'd23816; ROM4[5788]<=16'd57300;
ROM1[5789]<=16'd4857; ROM2[5789]<=16'd0; ROM3[5789]<=16'd23832; ROM4[5789]<=16'd57327;
ROM1[5790]<=16'd4880; ROM2[5790]<=16'd0; ROM3[5790]<=16'd23807; ROM4[5790]<=16'd57316;
ROM1[5791]<=16'd4858; ROM2[5791]<=16'd0; ROM3[5791]<=16'd23770; ROM4[5791]<=16'd57281;
ROM1[5792]<=16'd4842; ROM2[5792]<=16'd0; ROM3[5792]<=16'd23768; ROM4[5792]<=16'd57272;
ROM1[5793]<=16'd4830; ROM2[5793]<=16'd0; ROM3[5793]<=16'd23786; ROM4[5793]<=16'd57284;
ROM1[5794]<=16'd4834; ROM2[5794]<=16'd0; ROM3[5794]<=16'd23813; ROM4[5794]<=16'd57306;
ROM1[5795]<=16'd4835; ROM2[5795]<=16'd0; ROM3[5795]<=16'd23833; ROM4[5795]<=16'd57323;
ROM1[5796]<=16'd4829; ROM2[5796]<=16'd0; ROM3[5796]<=16'd23832; ROM4[5796]<=16'd57320;
ROM1[5797]<=16'd4828; ROM2[5797]<=16'd0; ROM3[5797]<=16'd23807; ROM4[5797]<=16'd57300;
ROM1[5798]<=16'd4853; ROM2[5798]<=16'd0; ROM3[5798]<=16'd23788; ROM4[5798]<=16'd57289;
ROM1[5799]<=16'd4877; ROM2[5799]<=16'd0; ROM3[5799]<=16'd23783; ROM4[5799]<=16'd57294;
ROM1[5800]<=16'd4864; ROM2[5800]<=16'd0; ROM3[5800]<=16'd23780; ROM4[5800]<=16'd57296;
ROM1[5801]<=16'd4837; ROM2[5801]<=16'd0; ROM3[5801]<=16'd23781; ROM4[5801]<=16'd57285;
ROM1[5802]<=16'd4823; ROM2[5802]<=16'd0; ROM3[5802]<=16'd23789; ROM4[5802]<=16'd57289;
ROM1[5803]<=16'd4819; ROM2[5803]<=16'd0; ROM3[5803]<=16'd23795; ROM4[5803]<=16'd57295;
ROM1[5804]<=16'd4800; ROM2[5804]<=16'd0; ROM3[5804]<=16'd23793; ROM4[5804]<=16'd57285;
ROM1[5805]<=16'd4805; ROM2[5805]<=16'd0; ROM3[5805]<=16'd23792; ROM4[5805]<=16'd57285;
ROM1[5806]<=16'd4822; ROM2[5806]<=16'd0; ROM3[5806]<=16'd23777; ROM4[5806]<=16'd57278;
ROM1[5807]<=16'd4845; ROM2[5807]<=16'd0; ROM3[5807]<=16'd23770; ROM4[5807]<=16'd57281;
ROM1[5808]<=16'd4842; ROM2[5808]<=16'd0; ROM3[5808]<=16'd23770; ROM4[5808]<=16'd57281;
ROM1[5809]<=16'd4816; ROM2[5809]<=16'd0; ROM3[5809]<=16'd23765; ROM4[5809]<=16'd57274;
ROM1[5810]<=16'd4799; ROM2[5810]<=16'd0; ROM3[5810]<=16'd23769; ROM4[5810]<=16'd57272;
ROM1[5811]<=16'd4789; ROM2[5811]<=16'd0; ROM3[5811]<=16'd23773; ROM4[5811]<=16'd57269;
ROM1[5812]<=16'd4777; ROM2[5812]<=16'd0; ROM3[5812]<=16'd23774; ROM4[5812]<=16'd57274;
ROM1[5813]<=16'd4778; ROM2[5813]<=16'd0; ROM3[5813]<=16'd23776; ROM4[5813]<=16'd57274;
ROM1[5814]<=16'd4800; ROM2[5814]<=16'd0; ROM3[5814]<=16'd23771; ROM4[5814]<=16'd57274;
ROM1[5815]<=16'd4826; ROM2[5815]<=16'd0; ROM3[5815]<=16'd23750; ROM4[5815]<=16'd57268;
ROM1[5816]<=16'd4837; ROM2[5816]<=16'd0; ROM3[5816]<=16'd23740; ROM4[5816]<=16'd57261;
ROM1[5817]<=16'd4825; ROM2[5817]<=16'd0; ROM3[5817]<=16'd23746; ROM4[5817]<=16'd57263;
ROM1[5818]<=16'd4809; ROM2[5818]<=16'd0; ROM3[5818]<=16'd23758; ROM4[5818]<=16'd57270;
ROM1[5819]<=16'd4801; ROM2[5819]<=16'd0; ROM3[5819]<=16'd23773; ROM4[5819]<=16'd57276;
ROM1[5820]<=16'd4771; ROM2[5820]<=16'd0; ROM3[5820]<=16'd23761; ROM4[5820]<=16'd57263;
ROM1[5821]<=16'd4762; ROM2[5821]<=16'd0; ROM3[5821]<=16'd23758; ROM4[5821]<=16'd57261;
ROM1[5822]<=16'd4779; ROM2[5822]<=16'd0; ROM3[5822]<=16'd23757; ROM4[5822]<=16'd57264;
ROM1[5823]<=16'd4809; ROM2[5823]<=16'd0; ROM3[5823]<=16'd23739; ROM4[5823]<=16'd57258;
ROM1[5824]<=16'd4838; ROM2[5824]<=16'd0; ROM3[5824]<=16'd23743; ROM4[5824]<=16'd57266;
ROM1[5825]<=16'd4833; ROM2[5825]<=16'd0; ROM3[5825]<=16'd23755; ROM4[5825]<=16'd57271;
ROM1[5826]<=16'd4819; ROM2[5826]<=16'd0; ROM3[5826]<=16'd23770; ROM4[5826]<=16'd57277;
ROM1[5827]<=16'd4809; ROM2[5827]<=16'd0; ROM3[5827]<=16'd23785; ROM4[5827]<=16'd57283;
ROM1[5828]<=16'd4806; ROM2[5828]<=16'd0; ROM3[5828]<=16'd23799; ROM4[5828]<=16'd57293;
ROM1[5829]<=16'd4805; ROM2[5829]<=16'd0; ROM3[5829]<=16'd23804; ROM4[5829]<=16'd57296;
ROM1[5830]<=16'd4809; ROM2[5830]<=16'd0; ROM3[5830]<=16'd23798; ROM4[5830]<=16'd57292;
ROM1[5831]<=16'd4837; ROM2[5831]<=16'd0; ROM3[5831]<=16'd23794; ROM4[5831]<=16'd57295;
ROM1[5832]<=16'd4873; ROM2[5832]<=16'd0; ROM3[5832]<=16'd23788; ROM4[5832]<=16'd57299;
ROM1[5833]<=16'd4863; ROM2[5833]<=16'd0; ROM3[5833]<=16'd23775; ROM4[5833]<=16'd57289;
ROM1[5834]<=16'd4839; ROM2[5834]<=16'd0; ROM3[5834]<=16'd23774; ROM4[5834]<=16'd57285;
ROM1[5835]<=16'd4822; ROM2[5835]<=16'd0; ROM3[5835]<=16'd23786; ROM4[5835]<=16'd57290;
ROM1[5836]<=16'd4808; ROM2[5836]<=16'd0; ROM3[5836]<=16'd23790; ROM4[5836]<=16'd57291;
ROM1[5837]<=16'd4802; ROM2[5837]<=16'd0; ROM3[5837]<=16'd23799; ROM4[5837]<=16'd57293;
ROM1[5838]<=16'd4808; ROM2[5838]<=16'd0; ROM3[5838]<=16'd23799; ROM4[5838]<=16'd57292;
ROM1[5839]<=16'd4816; ROM2[5839]<=16'd0; ROM3[5839]<=16'd23774; ROM4[5839]<=16'd57279;
ROM1[5840]<=16'd4844; ROM2[5840]<=16'd0; ROM3[5840]<=16'd23762; ROM4[5840]<=16'd57273;
ROM1[5841]<=16'd4880; ROM2[5841]<=16'd0; ROM3[5841]<=16'd23785; ROM4[5841]<=16'd57300;
ROM1[5842]<=16'd4874; ROM2[5842]<=16'd0; ROM3[5842]<=16'd23797; ROM4[5842]<=16'd57311;
ROM1[5843]<=16'd4842; ROM2[5843]<=16'd0; ROM3[5843]<=16'd23795; ROM4[5843]<=16'd57300;
ROM1[5844]<=16'd4810; ROM2[5844]<=16'd0; ROM3[5844]<=16'd23786; ROM4[5844]<=16'd57280;
ROM1[5845]<=16'd4768; ROM2[5845]<=16'd0; ROM3[5845]<=16'd23769; ROM4[5845]<=16'd57252;
ROM1[5846]<=16'd4759; ROM2[5846]<=16'd0; ROM3[5846]<=16'd23768; ROM4[5846]<=16'd57245;
ROM1[5847]<=16'd4789; ROM2[5847]<=16'd0; ROM3[5847]<=16'd23777; ROM4[5847]<=16'd57257;
ROM1[5848]<=16'd4827; ROM2[5848]<=16'd0; ROM3[5848]<=16'd23773; ROM4[5848]<=16'd57263;
ROM1[5849]<=16'd4851; ROM2[5849]<=16'd0; ROM3[5849]<=16'd23762; ROM4[5849]<=16'd57265;
ROM1[5850]<=16'd4842; ROM2[5850]<=16'd0; ROM3[5850]<=16'd23760; ROM4[5850]<=16'd57264;
ROM1[5851]<=16'd4823; ROM2[5851]<=16'd0; ROM3[5851]<=16'd23765; ROM4[5851]<=16'd57259;
ROM1[5852]<=16'd4809; ROM2[5852]<=16'd0; ROM3[5852]<=16'd23771; ROM4[5852]<=16'd57256;
ROM1[5853]<=16'd4795; ROM2[5853]<=16'd0; ROM3[5853]<=16'd23781; ROM4[5853]<=16'd57263;
ROM1[5854]<=16'd4779; ROM2[5854]<=16'd0; ROM3[5854]<=16'd23782; ROM4[5854]<=16'd57261;
ROM1[5855]<=16'd4785; ROM2[5855]<=16'd0; ROM3[5855]<=16'd23773; ROM4[5855]<=16'd57259;
ROM1[5856]<=16'd4822; ROM2[5856]<=16'd0; ROM3[5856]<=16'd23765; ROM4[5856]<=16'd57263;
ROM1[5857]<=16'd4855; ROM2[5857]<=16'd0; ROM3[5857]<=16'd23750; ROM4[5857]<=16'd57262;
ROM1[5858]<=16'd4844; ROM2[5858]<=16'd0; ROM3[5858]<=16'd23741; ROM4[5858]<=16'd57254;
ROM1[5859]<=16'd4823; ROM2[5859]<=16'd0; ROM3[5859]<=16'd23745; ROM4[5859]<=16'd57251;
ROM1[5860]<=16'd4810; ROM2[5860]<=16'd0; ROM3[5860]<=16'd23753; ROM4[5860]<=16'd57256;
ROM1[5861]<=16'd4813; ROM2[5861]<=16'd0; ROM3[5861]<=16'd23763; ROM4[5861]<=16'd57261;
ROM1[5862]<=16'd4811; ROM2[5862]<=16'd0; ROM3[5862]<=16'd23774; ROM4[5862]<=16'd57265;
ROM1[5863]<=16'd4824; ROM2[5863]<=16'd0; ROM3[5863]<=16'd23787; ROM4[5863]<=16'd57277;
ROM1[5864]<=16'd4859; ROM2[5864]<=16'd0; ROM3[5864]<=16'd23796; ROM4[5864]<=16'd57294;
ROM1[5865]<=16'd4882; ROM2[5865]<=16'd0; ROM3[5865]<=16'd23777; ROM4[5865]<=16'd57289;
ROM1[5866]<=16'd4892; ROM2[5866]<=16'd0; ROM3[5866]<=16'd23765; ROM4[5866]<=16'd57281;
ROM1[5867]<=16'd4889; ROM2[5867]<=16'd0; ROM3[5867]<=16'd23771; ROM4[5867]<=16'd57284;
ROM1[5868]<=16'd4859; ROM2[5868]<=16'd0; ROM3[5868]<=16'd23776; ROM4[5868]<=16'd57281;
ROM1[5869]<=16'd4863; ROM2[5869]<=16'd0; ROM3[5869]<=16'd23799; ROM4[5869]<=16'd57295;
ROM1[5870]<=16'd4880; ROM2[5870]<=16'd0; ROM3[5870]<=16'd23816; ROM4[5870]<=16'd57310;
ROM1[5871]<=16'd4880; ROM2[5871]<=16'd0; ROM3[5871]<=16'd23801; ROM4[5871]<=16'd57297;
ROM1[5872]<=16'd4904; ROM2[5872]<=16'd0; ROM3[5872]<=16'd23782; ROM4[5872]<=16'd57289;
ROM1[5873]<=16'd4944; ROM2[5873]<=16'd0; ROM3[5873]<=16'd23767; ROM4[5873]<=16'd57290;
ROM1[5874]<=16'd4994; ROM2[5874]<=16'd0; ROM3[5874]<=16'd23777; ROM4[5874]<=16'd57311;
ROM1[5875]<=16'd5019; ROM2[5875]<=16'd0; ROM3[5875]<=16'd23804; ROM4[5875]<=16'd57339;
ROM1[5876]<=16'd5011; ROM2[5876]<=16'd0; ROM3[5876]<=16'd23811; ROM4[5876]<=16'd57344;
ROM1[5877]<=16'd5002; ROM2[5877]<=16'd0; ROM3[5877]<=16'd23808; ROM4[5877]<=16'd57337;
ROM1[5878]<=16'd5002; ROM2[5878]<=16'd0; ROM3[5878]<=16'd23812; ROM4[5878]<=16'd57338;
ROM1[5879]<=16'd5013; ROM2[5879]<=16'd0; ROM3[5879]<=16'd23819; ROM4[5879]<=16'd57344;
ROM1[5880]<=16'd5054; ROM2[5880]<=16'd0; ROM3[5880]<=16'd23837; ROM4[5880]<=16'd57364;
ROM1[5881]<=16'd5089; ROM2[5881]<=16'd0; ROM3[5881]<=16'd23830; ROM4[5881]<=16'd57366;
ROM1[5882]<=16'd5107; ROM2[5882]<=16'd0; ROM3[5882]<=16'd23799; ROM4[5882]<=16'd57348;
ROM1[5883]<=16'd5117; ROM2[5883]<=16'd0; ROM3[5883]<=16'd23800; ROM4[5883]<=16'd57350;
ROM1[5884]<=16'd5114; ROM2[5884]<=16'd0; ROM3[5884]<=16'd23809; ROM4[5884]<=16'd57351;
ROM1[5885]<=16'd5108; ROM2[5885]<=16'd0; ROM3[5885]<=16'd23819; ROM4[5885]<=16'd57352;
ROM1[5886]<=16'd5108; ROM2[5886]<=16'd0; ROM3[5886]<=16'd23830; ROM4[5886]<=16'd57359;
ROM1[5887]<=16'd5104; ROM2[5887]<=16'd0; ROM3[5887]<=16'd23831; ROM4[5887]<=16'd57359;
ROM1[5888]<=16'd5116; ROM2[5888]<=16'd0; ROM3[5888]<=16'd23827; ROM4[5888]<=16'd57365;
ROM1[5889]<=16'd5156; ROM2[5889]<=16'd0; ROM3[5889]<=16'd23829; ROM4[5889]<=16'd57376;
ROM1[5890]<=16'd5200; ROM2[5890]<=16'd0; ROM3[5890]<=16'd23825; ROM4[5890]<=16'd57382;
ROM1[5891]<=16'd5217; ROM2[5891]<=16'd0; ROM3[5891]<=16'd23828; ROM4[5891]<=16'd57390;
ROM1[5892]<=16'd5211; ROM2[5892]<=16'd0; ROM3[5892]<=16'd23839; ROM4[5892]<=16'd57398;
ROM1[5893]<=16'd5193; ROM2[5893]<=16'd0; ROM3[5893]<=16'd23845; ROM4[5893]<=16'd57396;
ROM1[5894]<=16'd5167; ROM2[5894]<=16'd0; ROM3[5894]<=16'd23837; ROM4[5894]<=16'd57383;
ROM1[5895]<=16'd5144; ROM2[5895]<=16'd0; ROM3[5895]<=16'd23829; ROM4[5895]<=16'd57368;
ROM1[5896]<=16'd5143; ROM2[5896]<=16'd0; ROM3[5896]<=16'd23829; ROM4[5896]<=16'd57367;
ROM1[5897]<=16'd5173; ROM2[5897]<=16'd0; ROM3[5897]<=16'd23835; ROM4[5897]<=16'd57381;
ROM1[5898]<=16'd5213; ROM2[5898]<=16'd0; ROM3[5898]<=16'd23840; ROM4[5898]<=16'd57394;
ROM1[5899]<=16'd5230; ROM2[5899]<=16'd0; ROM3[5899]<=16'd23837; ROM4[5899]<=16'd57395;
ROM1[5900]<=16'd5209; ROM2[5900]<=16'd0; ROM3[5900]<=16'd23833; ROM4[5900]<=16'd57384;
ROM1[5901]<=16'd5172; ROM2[5901]<=16'd0; ROM3[5901]<=16'd23829; ROM4[5901]<=16'd57372;
ROM1[5902]<=16'd5148; ROM2[5902]<=16'd0; ROM3[5902]<=16'd23831; ROM4[5902]<=16'd57369;
ROM1[5903]<=16'd5134; ROM2[5903]<=16'd0; ROM3[5903]<=16'd23839; ROM4[5903]<=16'd57371;
ROM1[5904]<=16'd5114; ROM2[5904]<=16'd0; ROM3[5904]<=16'd23840; ROM4[5904]<=16'd57365;
ROM1[5905]<=16'd5109; ROM2[5905]<=16'd0; ROM3[5905]<=16'd23832; ROM4[5905]<=16'd57357;
ROM1[5906]<=16'd5135; ROM2[5906]<=16'd0; ROM3[5906]<=16'd23824; ROM4[5906]<=16'd57360;
ROM1[5907]<=16'd5158; ROM2[5907]<=16'd0; ROM3[5907]<=16'd23809; ROM4[5907]<=16'd57358;
ROM1[5908]<=16'd5150; ROM2[5908]<=16'd0; ROM3[5908]<=16'd23804; ROM4[5908]<=16'd57357;
ROM1[5909]<=16'd5123; ROM2[5909]<=16'd0; ROM3[5909]<=16'd23808; ROM4[5909]<=16'd57354;
ROM1[5910]<=16'd5101; ROM2[5910]<=16'd0; ROM3[5910]<=16'd23812; ROM4[5910]<=16'd57347;
ROM1[5911]<=16'd5103; ROM2[5911]<=16'd0; ROM3[5911]<=16'd23835; ROM4[5911]<=16'd57368;
ROM1[5912]<=16'd5104; ROM2[5912]<=16'd0; ROM3[5912]<=16'd23860; ROM4[5912]<=16'd57388;
ROM1[5913]<=16'd5059; ROM2[5913]<=16'd0; ROM3[5913]<=16'd23822; ROM4[5913]<=16'd57350;
ROM1[5914]<=16'd5034; ROM2[5914]<=16'd0; ROM3[5914]<=16'd23780; ROM4[5914]<=16'd57321;
ROM1[5915]<=16'd5069; ROM2[5915]<=16'd0; ROM3[5915]<=16'd23772; ROM4[5915]<=16'd57325;
ROM1[5916]<=16'd5074; ROM2[5916]<=16'd0; ROM3[5916]<=16'd23763; ROM4[5916]<=16'd57318;
ROM1[5917]<=16'd5081; ROM2[5917]<=16'd0; ROM3[5917]<=16'd23791; ROM4[5917]<=16'd57340;
ROM1[5918]<=16'd5074; ROM2[5918]<=16'd0; ROM3[5918]<=16'd23817; ROM4[5918]<=16'd57360;
ROM1[5919]<=16'd5020; ROM2[5919]<=16'd0; ROM3[5919]<=16'd23797; ROM4[5919]<=16'd57330;
ROM1[5920]<=16'd4988; ROM2[5920]<=16'd0; ROM3[5920]<=16'd23791; ROM4[5920]<=16'd57316;
ROM1[5921]<=16'd5009; ROM2[5921]<=16'd0; ROM3[5921]<=16'd23817; ROM4[5921]<=16'd57342;
ROM1[5922]<=16'd5021; ROM2[5922]<=16'd0; ROM3[5922]<=16'd23812; ROM4[5922]<=16'd57338;
ROM1[5923]<=16'd5026; ROM2[5923]<=16'd0; ROM3[5923]<=16'd23785; ROM4[5923]<=16'd57320;
ROM1[5924]<=16'd5030; ROM2[5924]<=16'd0; ROM3[5924]<=16'd23774; ROM4[5924]<=16'd57315;
ROM1[5925]<=16'd5014; ROM2[5925]<=16'd0; ROM3[5925]<=16'd23775; ROM4[5925]<=16'd57313;
ROM1[5926]<=16'd5008; ROM2[5926]<=16'd0; ROM3[5926]<=16'd23798; ROM4[5926]<=16'd57331;
ROM1[5927]<=16'd4998; ROM2[5927]<=16'd0; ROM3[5927]<=16'd23819; ROM4[5927]<=16'd57341;
ROM1[5928]<=16'd4973; ROM2[5928]<=16'd0; ROM3[5928]<=16'd23821; ROM4[5928]<=16'd57332;
ROM1[5929]<=16'd4954; ROM2[5929]<=16'd0; ROM3[5929]<=16'd23820; ROM4[5929]<=16'd57328;
ROM1[5930]<=16'd4965; ROM2[5930]<=16'd0; ROM3[5930]<=16'd23831; ROM4[5930]<=16'd57334;
ROM1[5931]<=16'd5003; ROM2[5931]<=16'd0; ROM3[5931]<=16'd23836; ROM4[5931]<=16'd57351;
ROM1[5932]<=16'd5012; ROM2[5932]<=16'd0; ROM3[5932]<=16'd23810; ROM4[5932]<=16'd57338;
ROM1[5933]<=16'd4995; ROM2[5933]<=16'd0; ROM3[5933]<=16'd23798; ROM4[5933]<=16'd57324;
ROM1[5934]<=16'd4972; ROM2[5934]<=16'd0; ROM3[5934]<=16'd23800; ROM4[5934]<=16'd57318;
ROM1[5935]<=16'd4946; ROM2[5935]<=16'd0; ROM3[5935]<=16'd23801; ROM4[5935]<=16'd57312;
ROM1[5936]<=16'd4940; ROM2[5936]<=16'd0; ROM3[5936]<=16'd23817; ROM4[5936]<=16'd57325;
ROM1[5937]<=16'd4924; ROM2[5937]<=16'd0; ROM3[5937]<=16'd23823; ROM4[5937]<=16'd57326;
ROM1[5938]<=16'd4906; ROM2[5938]<=16'd0; ROM3[5938]<=16'd23806; ROM4[5938]<=16'd57308;
ROM1[5939]<=16'd4909; ROM2[5939]<=16'd0; ROM3[5939]<=16'd23786; ROM4[5939]<=16'd57298;
ROM1[5940]<=16'd4946; ROM2[5940]<=16'd0; ROM3[5940]<=16'd23779; ROM4[5940]<=16'd57304;
ROM1[5941]<=16'd4965; ROM2[5941]<=16'd0; ROM3[5941]<=16'd23785; ROM4[5941]<=16'd57313;
ROM1[5942]<=16'd4965; ROM2[5942]<=16'd0; ROM3[5942]<=16'd23799; ROM4[5942]<=16'd57326;
ROM1[5943]<=16'd4933; ROM2[5943]<=16'd0; ROM3[5943]<=16'd23791; ROM4[5943]<=16'd57309;
ROM1[5944]<=16'd4897; ROM2[5944]<=16'd0; ROM3[5944]<=16'd23778; ROM4[5944]<=16'd57289;
ROM1[5945]<=16'd4880; ROM2[5945]<=16'd0; ROM3[5945]<=16'd23782; ROM4[5945]<=16'd57290;
ROM1[5946]<=16'd4863; ROM2[5946]<=16'd0; ROM3[5946]<=16'd23780; ROM4[5946]<=16'd57279;
ROM1[5947]<=16'd4877; ROM2[5947]<=16'd0; ROM3[5947]<=16'd23781; ROM4[5947]<=16'd57281;
ROM1[5948]<=16'd4917; ROM2[5948]<=16'd0; ROM3[5948]<=16'd23777; ROM4[5948]<=16'd57291;
ROM1[5949]<=16'd4924; ROM2[5949]<=16'd0; ROM3[5949]<=16'd23758; ROM4[5949]<=16'd57281;
ROM1[5950]<=16'd4906; ROM2[5950]<=16'd0; ROM3[5950]<=16'd23749; ROM4[5950]<=16'd57274;
ROM1[5951]<=16'd4896; ROM2[5951]<=16'd0; ROM3[5951]<=16'd23765; ROM4[5951]<=16'd57285;
ROM1[5952]<=16'd4893; ROM2[5952]<=16'd0; ROM3[5952]<=16'd23791; ROM4[5952]<=16'd57304;
ROM1[5953]<=16'd4878; ROM2[5953]<=16'd0; ROM3[5953]<=16'd23796; ROM4[5953]<=16'd57303;
ROM1[5954]<=16'd4852; ROM2[5954]<=16'd0; ROM3[5954]<=16'd23782; ROM4[5954]<=16'd57285;
ROM1[5955]<=16'd4851; ROM2[5955]<=16'd0; ROM3[5955]<=16'd23774; ROM4[5955]<=16'd57279;
ROM1[5956]<=16'd4872; ROM2[5956]<=16'd0; ROM3[5956]<=16'd23760; ROM4[5956]<=16'd57270;
ROM1[5957]<=16'd4903; ROM2[5957]<=16'd0; ROM3[5957]<=16'd23751; ROM4[5957]<=16'd57270;
ROM1[5958]<=16'd4910; ROM2[5958]<=16'd0; ROM3[5958]<=16'd23754; ROM4[5958]<=16'd57276;
ROM1[5959]<=16'd4889; ROM2[5959]<=16'd0; ROM3[5959]<=16'd23749; ROM4[5959]<=16'd57272;
ROM1[5960]<=16'd4865; ROM2[5960]<=16'd0; ROM3[5960]<=16'd23749; ROM4[5960]<=16'd57263;
ROM1[5961]<=16'd4850; ROM2[5961]<=16'd0; ROM3[5961]<=16'd23756; ROM4[5961]<=16'd57262;
ROM1[5962]<=16'd4840; ROM2[5962]<=16'd0; ROM3[5962]<=16'd23765; ROM4[5962]<=16'd57267;
ROM1[5963]<=16'd4853; ROM2[5963]<=16'd0; ROM3[5963]<=16'd23775; ROM4[5963]<=16'd57275;
ROM1[5964]<=16'd4878; ROM2[5964]<=16'd0; ROM3[5964]<=16'd23770; ROM4[5964]<=16'd57277;
ROM1[5965]<=16'd4896; ROM2[5965]<=16'd0; ROM3[5965]<=16'd23742; ROM4[5965]<=16'd57263;
ROM1[5966]<=16'd4897; ROM2[5966]<=16'd0; ROM3[5966]<=16'd23735; ROM4[5966]<=16'd57256;
ROM1[5967]<=16'd4876; ROM2[5967]<=16'd0; ROM3[5967]<=16'd23736; ROM4[5967]<=16'd57250;
ROM1[5968]<=16'd4851; ROM2[5968]<=16'd0; ROM3[5968]<=16'd23737; ROM4[5968]<=16'd57246;
ROM1[5969]<=16'd4842; ROM2[5969]<=16'd0; ROM3[5969]<=16'd23752; ROM4[5969]<=16'd57254;
ROM1[5970]<=16'd4836; ROM2[5970]<=16'd0; ROM3[5970]<=16'd23776; ROM4[5970]<=16'd57270;
ROM1[5971]<=16'd4835; ROM2[5971]<=16'd0; ROM3[5971]<=16'd23776; ROM4[5971]<=16'd57270;
ROM1[5972]<=16'd4840; ROM2[5972]<=16'd0; ROM3[5972]<=16'd23762; ROM4[5972]<=16'd57261;
ROM1[5973]<=16'd4865; ROM2[5973]<=16'd0; ROM3[5973]<=16'd23750; ROM4[5973]<=16'd57259;
ROM1[5974]<=16'd4882; ROM2[5974]<=16'd0; ROM3[5974]<=16'd23734; ROM4[5974]<=16'd57253;
ROM1[5975]<=16'd4866; ROM2[5975]<=16'd0; ROM3[5975]<=16'd23739; ROM4[5975]<=16'd57251;
ROM1[5976]<=16'd4848; ROM2[5976]<=16'd0; ROM3[5976]<=16'd23746; ROM4[5976]<=16'd57247;
ROM1[5977]<=16'd4841; ROM2[5977]<=16'd0; ROM3[5977]<=16'd23756; ROM4[5977]<=16'd57248;
ROM1[5978]<=16'd4832; ROM2[5978]<=16'd0; ROM3[5978]<=16'd23766; ROM4[5978]<=16'd57259;
ROM1[5979]<=16'd4823; ROM2[5979]<=16'd0; ROM3[5979]<=16'd23769; ROM4[5979]<=16'd57260;
ROM1[5980]<=16'd4838; ROM2[5980]<=16'd0; ROM3[5980]<=16'd23772; ROM4[5980]<=16'd57264;
ROM1[5981]<=16'd4903; ROM2[5981]<=16'd0; ROM3[5981]<=16'd23797; ROM4[5981]<=16'd57302;
ROM1[5982]<=16'd4935; ROM2[5982]<=16'd0; ROM3[5982]<=16'd23786; ROM4[5982]<=16'd57301;
ROM1[5983]<=16'd4897; ROM2[5983]<=16'd0; ROM3[5983]<=16'd23750; ROM4[5983]<=16'd57267;
ROM1[5984]<=16'd4873; ROM2[5984]<=16'd0; ROM3[5984]<=16'd23754; ROM4[5984]<=16'd57262;
ROM1[5985]<=16'd4850; ROM2[5985]<=16'd0; ROM3[5985]<=16'd23759; ROM4[5985]<=16'd57259;
ROM1[5986]<=16'd4827; ROM2[5986]<=16'd0; ROM3[5986]<=16'd23754; ROM4[5986]<=16'd57251;
ROM1[5987]<=16'd4823; ROM2[5987]<=16'd0; ROM3[5987]<=16'd23767; ROM4[5987]<=16'd57258;
ROM1[5988]<=16'd4834; ROM2[5988]<=16'd0; ROM3[5988]<=16'd23777; ROM4[5988]<=16'd57271;
ROM1[5989]<=16'd4844; ROM2[5989]<=16'd0; ROM3[5989]<=16'd23759; ROM4[5989]<=16'd57263;
ROM1[5990]<=16'd4873; ROM2[5990]<=16'd0; ROM3[5990]<=16'd23741; ROM4[5990]<=16'd57261;
ROM1[5991]<=16'd4892; ROM2[5991]<=16'd0; ROM3[5991]<=16'd23744; ROM4[5991]<=16'd57274;
ROM1[5992]<=16'd4894; ROM2[5992]<=16'd0; ROM3[5992]<=16'd23766; ROM4[5992]<=16'd57290;
ROM1[5993]<=16'd4858; ROM2[5993]<=16'd0; ROM3[5993]<=16'd23756; ROM4[5993]<=16'd57277;
ROM1[5994]<=16'd4817; ROM2[5994]<=16'd0; ROM3[5994]<=16'd23737; ROM4[5994]<=16'd57254;
ROM1[5995]<=16'd4816; ROM2[5995]<=16'd0; ROM3[5995]<=16'd23760; ROM4[5995]<=16'd57269;
ROM1[5996]<=16'd4813; ROM2[5996]<=16'd0; ROM3[5996]<=16'd23763; ROM4[5996]<=16'd57271;
ROM1[5997]<=16'd4833; ROM2[5997]<=16'd0; ROM3[5997]<=16'd23758; ROM4[5997]<=16'd57274;
ROM1[5998]<=16'd4878; ROM2[5998]<=16'd0; ROM3[5998]<=16'd23766; ROM4[5998]<=16'd57283;
ROM1[5999]<=16'd4900; ROM2[5999]<=16'd0; ROM3[5999]<=16'd23761; ROM4[5999]<=16'd57285;
ROM1[6000]<=16'd4875; ROM2[6000]<=16'd0; ROM3[6000]<=16'd23753; ROM4[6000]<=16'd57276;
ROM1[6001]<=16'd4846; ROM2[6001]<=16'd0; ROM3[6001]<=16'd23755; ROM4[6001]<=16'd57270;
ROM1[6002]<=16'd4838; ROM2[6002]<=16'd0; ROM3[6002]<=16'd23776; ROM4[6002]<=16'd57282;
ROM1[6003]<=16'd4821; ROM2[6003]<=16'd0; ROM3[6003]<=16'd23789; ROM4[6003]<=16'd57282;
ROM1[6004]<=16'd4806; ROM2[6004]<=16'd0; ROM3[6004]<=16'd23784; ROM4[6004]<=16'd57276;
ROM1[6005]<=16'd4821; ROM2[6005]<=16'd0; ROM3[6005]<=16'd23786; ROM4[6005]<=16'd57280;
ROM1[6006]<=16'd4857; ROM2[6006]<=16'd0; ROM3[6006]<=16'd23783; ROM4[6006]<=16'd57286;
ROM1[6007]<=16'd4884; ROM2[6007]<=16'd0; ROM3[6007]<=16'd23768; ROM4[6007]<=16'd57289;
ROM1[6008]<=16'd4883; ROM2[6008]<=16'd0; ROM3[6008]<=16'd23765; ROM4[6008]<=16'd57289;
ROM1[6009]<=16'd4860; ROM2[6009]<=16'd0; ROM3[6009]<=16'd23764; ROM4[6009]<=16'd57285;
ROM1[6010]<=16'd4844; ROM2[6010]<=16'd0; ROM3[6010]<=16'd23771; ROM4[6010]<=16'd57290;
ROM1[6011]<=16'd4837; ROM2[6011]<=16'd0; ROM3[6011]<=16'd23779; ROM4[6011]<=16'd57293;
ROM1[6012]<=16'd4826; ROM2[6012]<=16'd0; ROM3[6012]<=16'd23785; ROM4[6012]<=16'd57294;
ROM1[6013]<=16'd4825; ROM2[6013]<=16'd0; ROM3[6013]<=16'd23786; ROM4[6013]<=16'd57292;
ROM1[6014]<=16'd4847; ROM2[6014]<=16'd0; ROM3[6014]<=16'd23781; ROM4[6014]<=16'd57291;
ROM1[6015]<=16'd4881; ROM2[6015]<=16'd0; ROM3[6015]<=16'd23775; ROM4[6015]<=16'd57296;
ROM1[6016]<=16'd4877; ROM2[6016]<=16'd0; ROM3[6016]<=16'd23762; ROM4[6016]<=16'd57285;
ROM1[6017]<=16'd4876; ROM2[6017]<=16'd0; ROM3[6017]<=16'd23779; ROM4[6017]<=16'd57292;
ROM1[6018]<=16'd4868; ROM2[6018]<=16'd0; ROM3[6018]<=16'd23796; ROM4[6018]<=16'd57300;
ROM1[6019]<=16'd4847; ROM2[6019]<=16'd0; ROM3[6019]<=16'd23797; ROM4[6019]<=16'd57291;
ROM1[6020]<=16'd4830; ROM2[6020]<=16'd0; ROM3[6020]<=16'd23801; ROM4[6020]<=16'd57289;
ROM1[6021]<=16'd4819; ROM2[6021]<=16'd0; ROM3[6021]<=16'd23795; ROM4[6021]<=16'd57280;
ROM1[6022]<=16'd4821; ROM2[6022]<=16'd0; ROM3[6022]<=16'd23780; ROM4[6022]<=16'd57263;
ROM1[6023]<=16'd4846; ROM2[6023]<=16'd0; ROM3[6023]<=16'd23767; ROM4[6023]<=16'd57263;
ROM1[6024]<=16'd4873; ROM2[6024]<=16'd0; ROM3[6024]<=16'd23772; ROM4[6024]<=16'd57272;
ROM1[6025]<=16'd4861; ROM2[6025]<=16'd0; ROM3[6025]<=16'd23775; ROM4[6025]<=16'd57269;
ROM1[6026]<=16'd4849; ROM2[6026]<=16'd0; ROM3[6026]<=16'd23788; ROM4[6026]<=16'd57282;
ROM1[6027]<=16'd4840; ROM2[6027]<=16'd0; ROM3[6027]<=16'd23803; ROM4[6027]<=16'd57284;
ROM1[6028]<=16'd4811; ROM2[6028]<=16'd0; ROM3[6028]<=16'd23790; ROM4[6028]<=16'd57265;
ROM1[6029]<=16'd4804; ROM2[6029]<=16'd0; ROM3[6029]<=16'd23791; ROM4[6029]<=16'd57266;
ROM1[6030]<=16'd4820; ROM2[6030]<=16'd0; ROM3[6030]<=16'd23793; ROM4[6030]<=16'd57270;
ROM1[6031]<=16'd4842; ROM2[6031]<=16'd0; ROM3[6031]<=16'd23774; ROM4[6031]<=16'd57264;
ROM1[6032]<=16'd4871; ROM2[6032]<=16'd0; ROM3[6032]<=16'd23765; ROM4[6032]<=16'd57270;
ROM1[6033]<=16'd4865; ROM2[6033]<=16'd0; ROM3[6033]<=16'd23765; ROM4[6033]<=16'd57269;
ROM1[6034]<=16'd4836; ROM2[6034]<=16'd0; ROM3[6034]<=16'd23763; ROM4[6034]<=16'd57260;
ROM1[6035]<=16'd4819; ROM2[6035]<=16'd0; ROM3[6035]<=16'd23768; ROM4[6035]<=16'd57257;
ROM1[6036]<=16'd4813; ROM2[6036]<=16'd0; ROM3[6036]<=16'd23777; ROM4[6036]<=16'd57265;
ROM1[6037]<=16'd4814; ROM2[6037]<=16'd0; ROM3[6037]<=16'd23793; ROM4[6037]<=16'd57280;
ROM1[6038]<=16'd4821; ROM2[6038]<=16'd0; ROM3[6038]<=16'd23798; ROM4[6038]<=16'd57287;
ROM1[6039]<=16'd4824; ROM2[6039]<=16'd0; ROM3[6039]<=16'd23777; ROM4[6039]<=16'd57273;
ROM1[6040]<=16'd4852; ROM2[6040]<=16'd0; ROM3[6040]<=16'd23761; ROM4[6040]<=16'd57266;
ROM1[6041]<=16'd4859; ROM2[6041]<=16'd0; ROM3[6041]<=16'd23760; ROM4[6041]<=16'd57269;
ROM1[6042]<=16'd4852; ROM2[6042]<=16'd0; ROM3[6042]<=16'd23770; ROM4[6042]<=16'd57275;
ROM1[6043]<=16'd4847; ROM2[6043]<=16'd0; ROM3[6043]<=16'd23792; ROM4[6043]<=16'd57293;
ROM1[6044]<=16'd4833; ROM2[6044]<=16'd0; ROM3[6044]<=16'd23806; ROM4[6044]<=16'd57298;
ROM1[6045]<=16'd4812; ROM2[6045]<=16'd0; ROM3[6045]<=16'd23812; ROM4[6045]<=16'd57294;
ROM1[6046]<=16'd4800; ROM2[6046]<=16'd0; ROM3[6046]<=16'd23812; ROM4[6046]<=16'd57294;
ROM1[6047]<=16'd4822; ROM2[6047]<=16'd0; ROM3[6047]<=16'd23813; ROM4[6047]<=16'd57298;
ROM1[6048]<=16'd4863; ROM2[6048]<=16'd0; ROM3[6048]<=16'd23812; ROM4[6048]<=16'd57305;
ROM1[6049]<=16'd4899; ROM2[6049]<=16'd0; ROM3[6049]<=16'd23824; ROM4[6049]<=16'd57324;
ROM1[6050]<=16'd4894; ROM2[6050]<=16'd0; ROM3[6050]<=16'd23832; ROM4[6050]<=16'd57326;
ROM1[6051]<=16'd4856; ROM2[6051]<=16'd0; ROM3[6051]<=16'd23816; ROM4[6051]<=16'd57306;
ROM1[6052]<=16'd4837; ROM2[6052]<=16'd0; ROM3[6052]<=16'd23818; ROM4[6052]<=16'd57306;
ROM1[6053]<=16'd4817; ROM2[6053]<=16'd0; ROM3[6053]<=16'd23819; ROM4[6053]<=16'd57301;
ROM1[6054]<=16'd4798; ROM2[6054]<=16'd0; ROM3[6054]<=16'd23812; ROM4[6054]<=16'd57292;
ROM1[6055]<=16'd4811; ROM2[6055]<=16'd0; ROM3[6055]<=16'd23812; ROM4[6055]<=16'd57297;
ROM1[6056]<=16'd4847; ROM2[6056]<=16'd0; ROM3[6056]<=16'd23809; ROM4[6056]<=16'd57301;
ROM1[6057]<=16'd4874; ROM2[6057]<=16'd0; ROM3[6057]<=16'd23797; ROM4[6057]<=16'd57303;
ROM1[6058]<=16'd4880; ROM2[6058]<=16'd0; ROM3[6058]<=16'd23800; ROM4[6058]<=16'd57310;
ROM1[6059]<=16'd4870; ROM2[6059]<=16'd0; ROM3[6059]<=16'd23814; ROM4[6059]<=16'd57316;
ROM1[6060]<=16'd4845; ROM2[6060]<=16'd0; ROM3[6060]<=16'd23813; ROM4[6060]<=16'd57310;
ROM1[6061]<=16'd4823; ROM2[6061]<=16'd0; ROM3[6061]<=16'd23802; ROM4[6061]<=16'd57303;
ROM1[6062]<=16'd4808; ROM2[6062]<=16'd0; ROM3[6062]<=16'd23800; ROM4[6062]<=16'd57302;
ROM1[6063]<=16'd4815; ROM2[6063]<=16'd0; ROM3[6063]<=16'd23803; ROM4[6063]<=16'd57306;
ROM1[6064]<=16'd4838; ROM2[6064]<=16'd0; ROM3[6064]<=16'd23796; ROM4[6064]<=16'd57305;
ROM1[6065]<=16'd4869; ROM2[6065]<=16'd0; ROM3[6065]<=16'd23776; ROM4[6065]<=16'd57297;
ROM1[6066]<=16'd4871; ROM2[6066]<=16'd0; ROM3[6066]<=16'd23766; ROM4[6066]<=16'd57289;
ROM1[6067]<=16'd4861; ROM2[6067]<=16'd0; ROM3[6067]<=16'd23778; ROM4[6067]<=16'd57294;
ROM1[6068]<=16'd4842; ROM2[6068]<=16'd0; ROM3[6068]<=16'd23788; ROM4[6068]<=16'd57294;
ROM1[6069]<=16'd4818; ROM2[6069]<=16'd0; ROM3[6069]<=16'd23788; ROM4[6069]<=16'd57284;
ROM1[6070]<=16'd4812; ROM2[6070]<=16'd0; ROM3[6070]<=16'd23801; ROM4[6070]<=16'd57290;
ROM1[6071]<=16'd4816; ROM2[6071]<=16'd0; ROM3[6071]<=16'd23810; ROM4[6071]<=16'd57296;
ROM1[6072]<=16'd4835; ROM2[6072]<=16'd0; ROM3[6072]<=16'd23812; ROM4[6072]<=16'd57304;
ROM1[6073]<=16'd4855; ROM2[6073]<=16'd0; ROM3[6073]<=16'd23796; ROM4[6073]<=16'd57296;
ROM1[6074]<=16'd4858; ROM2[6074]<=16'd0; ROM3[6074]<=16'd23783; ROM4[6074]<=16'd57284;
ROM1[6075]<=16'd4848; ROM2[6075]<=16'd0; ROM3[6075]<=16'd23790; ROM4[6075]<=16'd57285;
ROM1[6076]<=16'd4840; ROM2[6076]<=16'd0; ROM3[6076]<=16'd23808; ROM4[6076]<=16'd57293;
ROM1[6077]<=16'd4845; ROM2[6077]<=16'd0; ROM3[6077]<=16'd23832; ROM4[6077]<=16'd57310;
ROM1[6078]<=16'd4816; ROM2[6078]<=16'd0; ROM3[6078]<=16'd23823; ROM4[6078]<=16'd57296;
ROM1[6079]<=16'd4785; ROM2[6079]<=16'd0; ROM3[6079]<=16'd23806; ROM4[6079]<=16'd57276;
ROM1[6080]<=16'd4790; ROM2[6080]<=16'd0; ROM3[6080]<=16'd23801; ROM4[6080]<=16'd57274;
ROM1[6081]<=16'd4834; ROM2[6081]<=16'd0; ROM3[6081]<=16'd23810; ROM4[6081]<=16'd57290;
ROM1[6082]<=16'd4876; ROM2[6082]<=16'd0; ROM3[6082]<=16'd23811; ROM4[6082]<=16'd57302;
ROM1[6083]<=16'd4864; ROM2[6083]<=16'd0; ROM3[6083]<=16'd23793; ROM4[6083]<=16'd57291;
ROM1[6084]<=16'd4843; ROM2[6084]<=16'd0; ROM3[6084]<=16'd23788; ROM4[6084]<=16'd57282;
ROM1[6085]<=16'd4823; ROM2[6085]<=16'd0; ROM3[6085]<=16'd23792; ROM4[6085]<=16'd57277;
ROM1[6086]<=16'd4813; ROM2[6086]<=16'd0; ROM3[6086]<=16'd23796; ROM4[6086]<=16'd57279;
ROM1[6087]<=16'd4814; ROM2[6087]<=16'd0; ROM3[6087]<=16'd23817; ROM4[6087]<=16'd57293;
ROM1[6088]<=16'd4805; ROM2[6088]<=16'd0; ROM3[6088]<=16'd23808; ROM4[6088]<=16'd57281;
ROM1[6089]<=16'd4804; ROM2[6089]<=16'd0; ROM3[6089]<=16'd23775; ROM4[6089]<=16'd57261;
ROM1[6090]<=16'd4850; ROM2[6090]<=16'd0; ROM3[6090]<=16'd23784; ROM4[6090]<=16'd57279;
ROM1[6091]<=16'd4874; ROM2[6091]<=16'd0; ROM3[6091]<=16'd23799; ROM4[6091]<=16'd57295;
ROM1[6092]<=16'd4860; ROM2[6092]<=16'd0; ROM3[6092]<=16'd23803; ROM4[6092]<=16'd57296;
ROM1[6093]<=16'd4839; ROM2[6093]<=16'd0; ROM3[6093]<=16'd23809; ROM4[6093]<=16'd57295;
ROM1[6094]<=16'd4821; ROM2[6094]<=16'd0; ROM3[6094]<=16'd23809; ROM4[6094]<=16'd57291;
ROM1[6095]<=16'd4803; ROM2[6095]<=16'd0; ROM3[6095]<=16'd23812; ROM4[6095]<=16'd57288;
ROM1[6096]<=16'd4798; ROM2[6096]<=16'd0; ROM3[6096]<=16'd23812; ROM4[6096]<=16'd57286;
ROM1[6097]<=16'd4821; ROM2[6097]<=16'd0; ROM3[6097]<=16'd23809; ROM4[6097]<=16'd57291;
ROM1[6098]<=16'd4847; ROM2[6098]<=16'd0; ROM3[6098]<=16'd23789; ROM4[6098]<=16'd57280;
ROM1[6099]<=16'd4856; ROM2[6099]<=16'd0; ROM3[6099]<=16'd23763; ROM4[6099]<=16'd57267;
ROM1[6100]<=16'd4845; ROM2[6100]<=16'd0; ROM3[6100]<=16'd23761; ROM4[6100]<=16'd57268;
ROM1[6101]<=16'd4818; ROM2[6101]<=16'd0; ROM3[6101]<=16'd23762; ROM4[6101]<=16'd57263;
ROM1[6102]<=16'd4806; ROM2[6102]<=16'd0; ROM3[6102]<=16'd23768; ROM4[6102]<=16'd57267;
ROM1[6103]<=16'd4818; ROM2[6103]<=16'd0; ROM3[6103]<=16'd23796; ROM4[6103]<=16'd57292;
ROM1[6104]<=16'd4813; ROM2[6104]<=16'd0; ROM3[6104]<=16'd23800; ROM4[6104]<=16'd57291;
ROM1[6105]<=16'd4807; ROM2[6105]<=16'd0; ROM3[6105]<=16'd23785; ROM4[6105]<=16'd57277;
ROM1[6106]<=16'd4824; ROM2[6106]<=16'd0; ROM3[6106]<=16'd23774; ROM4[6106]<=16'd57271;
ROM1[6107]<=16'd4848; ROM2[6107]<=16'd0; ROM3[6107]<=16'd23766; ROM4[6107]<=16'd57269;
ROM1[6108]<=16'd4855; ROM2[6108]<=16'd0; ROM3[6108]<=16'd23772; ROM4[6108]<=16'd57277;
ROM1[6109]<=16'd4851; ROM2[6109]<=16'd0; ROM3[6109]<=16'd23794; ROM4[6109]<=16'd57294;
ROM1[6110]<=16'd4846; ROM2[6110]<=16'd0; ROM3[6110]<=16'd23811; ROM4[6110]<=16'd57303;
ROM1[6111]<=16'd4822; ROM2[6111]<=16'd0; ROM3[6111]<=16'd23808; ROM4[6111]<=16'd57295;
ROM1[6112]<=16'd4800; ROM2[6112]<=16'd0; ROM3[6112]<=16'd23807; ROM4[6112]<=16'd57287;
ROM1[6113]<=16'd4803; ROM2[6113]<=16'd0; ROM3[6113]<=16'd23808; ROM4[6113]<=16'd57283;
ROM1[6114]<=16'd4820; ROM2[6114]<=16'd0; ROM3[6114]<=16'd23795; ROM4[6114]<=16'd57280;
ROM1[6115]<=16'd4861; ROM2[6115]<=16'd0; ROM3[6115]<=16'd23792; ROM4[6115]<=16'd57294;
ROM1[6116]<=16'd4872; ROM2[6116]<=16'd0; ROM3[6116]<=16'd23790; ROM4[6116]<=16'd57297;
ROM1[6117]<=16'd4851; ROM2[6117]<=16'd0; ROM3[6117]<=16'd23790; ROM4[6117]<=16'd57293;
ROM1[6118]<=16'd4840; ROM2[6118]<=16'd0; ROM3[6118]<=16'd23805; ROM4[6118]<=16'd57298;
ROM1[6119]<=16'd4829; ROM2[6119]<=16'd0; ROM3[6119]<=16'd23812; ROM4[6119]<=16'd57295;
ROM1[6120]<=16'd4825; ROM2[6120]<=16'd0; ROM3[6120]<=16'd23829; ROM4[6120]<=16'd57309;
ROM1[6121]<=16'd4813; ROM2[6121]<=16'd0; ROM3[6121]<=16'd23822; ROM4[6121]<=16'd57301;
ROM1[6122]<=16'd4805; ROM2[6122]<=16'd0; ROM3[6122]<=16'd23789; ROM4[6122]<=16'd57272;
ROM1[6123]<=16'd4831; ROM2[6123]<=16'd0; ROM3[6123]<=16'd23773; ROM4[6123]<=16'd57271;
ROM1[6124]<=16'd4848; ROM2[6124]<=16'd0; ROM3[6124]<=16'd23765; ROM4[6124]<=16'd57269;
ROM1[6125]<=16'd4846; ROM2[6125]<=16'd0; ROM3[6125]<=16'd23772; ROM4[6125]<=16'd57271;
ROM1[6126]<=16'd4834; ROM2[6126]<=16'd0; ROM3[6126]<=16'd23784; ROM4[6126]<=16'd57276;
ROM1[6127]<=16'd4814; ROM2[6127]<=16'd0; ROM3[6127]<=16'd23782; ROM4[6127]<=16'd57270;
ROM1[6128]<=16'd4793; ROM2[6128]<=16'd0; ROM3[6128]<=16'd23774; ROM4[6128]<=16'd57263;
ROM1[6129]<=16'd4793; ROM2[6129]<=16'd0; ROM3[6129]<=16'd23779; ROM4[6129]<=16'd57268;
ROM1[6130]<=16'd4811; ROM2[6130]<=16'd0; ROM3[6130]<=16'd23782; ROM4[6130]<=16'd57278;
ROM1[6131]<=16'd4837; ROM2[6131]<=16'd0; ROM3[6131]<=16'd23769; ROM4[6131]<=16'd57275;
ROM1[6132]<=16'd4864; ROM2[6132]<=16'd0; ROM3[6132]<=16'd23757; ROM4[6132]<=16'd57269;
ROM1[6133]<=16'd4855; ROM2[6133]<=16'd0; ROM3[6133]<=16'd23749; ROM4[6133]<=16'd57267;
ROM1[6134]<=16'd4856; ROM2[6134]<=16'd0; ROM3[6134]<=16'd23771; ROM4[6134]<=16'd57286;
ROM1[6135]<=16'd4848; ROM2[6135]<=16'd0; ROM3[6135]<=16'd23787; ROM4[6135]<=16'd57296;
ROM1[6136]<=16'd4819; ROM2[6136]<=16'd0; ROM3[6136]<=16'd23771; ROM4[6136]<=16'd57281;
ROM1[6137]<=16'd4815; ROM2[6137]<=16'd0; ROM3[6137]<=16'd23782; ROM4[6137]<=16'd57288;
ROM1[6138]<=16'd4813; ROM2[6138]<=16'd0; ROM3[6138]<=16'd23783; ROM4[6138]<=16'd57289;
ROM1[6139]<=16'd4813; ROM2[6139]<=16'd0; ROM3[6139]<=16'd23754; ROM4[6139]<=16'd57267;
ROM1[6140]<=16'd4843; ROM2[6140]<=16'd0; ROM3[6140]<=16'd23744; ROM4[6140]<=16'd57261;
ROM1[6141]<=16'd4854; ROM2[6141]<=16'd0; ROM3[6141]<=16'd23744; ROM4[6141]<=16'd57261;
ROM1[6142]<=16'd4837; ROM2[6142]<=16'd0; ROM3[6142]<=16'd23745; ROM4[6142]<=16'd57259;
ROM1[6143]<=16'd4823; ROM2[6143]<=16'd0; ROM3[6143]<=16'd23757; ROM4[6143]<=16'd57263;
ROM1[6144]<=16'd4813; ROM2[6144]<=16'd0; ROM3[6144]<=16'd23767; ROM4[6144]<=16'd57269;
ROM1[6145]<=16'd4799; ROM2[6145]<=16'd0; ROM3[6145]<=16'd23777; ROM4[6145]<=16'd57274;
ROM1[6146]<=16'd4803; ROM2[6146]<=16'd0; ROM3[6146]<=16'd23784; ROM4[6146]<=16'd57279;
ROM1[6147]<=16'd4829; ROM2[6147]<=16'd0; ROM3[6147]<=16'd23786; ROM4[6147]<=16'd57284;
ROM1[6148]<=16'd4852; ROM2[6148]<=16'd0; ROM3[6148]<=16'd23773; ROM4[6148]<=16'd57278;
ROM1[6149]<=16'd4854; ROM2[6149]<=16'd0; ROM3[6149]<=16'd23752; ROM4[6149]<=16'd57263;
ROM1[6150]<=16'd4832; ROM2[6150]<=16'd0; ROM3[6150]<=16'd23750; ROM4[6150]<=16'd57254;
ROM1[6151]<=16'd4815; ROM2[6151]<=16'd0; ROM3[6151]<=16'd23762; ROM4[6151]<=16'd57256;
ROM1[6152]<=16'd4817; ROM2[6152]<=16'd0; ROM3[6152]<=16'd23786; ROM4[6152]<=16'd57273;
ROM1[6153]<=16'd4811; ROM2[6153]<=16'd0; ROM3[6153]<=16'd23799; ROM4[6153]<=16'd57283;
ROM1[6154]<=16'd4803; ROM2[6154]<=16'd0; ROM3[6154]<=16'd23801; ROM4[6154]<=16'd57281;
ROM1[6155]<=16'd4811; ROM2[6155]<=16'd0; ROM3[6155]<=16'd23801; ROM4[6155]<=16'd57284;
ROM1[6156]<=16'd4837; ROM2[6156]<=16'd0; ROM3[6156]<=16'd23789; ROM4[6156]<=16'd57282;
ROM1[6157]<=16'd4879; ROM2[6157]<=16'd0; ROM3[6157]<=16'd23791; ROM4[6157]<=16'd57298;
ROM1[6158]<=16'd4876; ROM2[6158]<=16'd0; ROM3[6158]<=16'd23785; ROM4[6158]<=16'd57292;
ROM1[6159]<=16'd4839; ROM2[6159]<=16'd0; ROM3[6159]<=16'd23767; ROM4[6159]<=16'd57270;
ROM1[6160]<=16'd4828; ROM2[6160]<=16'd0; ROM3[6160]<=16'd23780; ROM4[6160]<=16'd57279;
ROM1[6161]<=16'd4821; ROM2[6161]<=16'd0; ROM3[6161]<=16'd23792; ROM4[6161]<=16'd57285;
ROM1[6162]<=16'd4809; ROM2[6162]<=16'd0; ROM3[6162]<=16'd23798; ROM4[6162]<=16'd57290;
ROM1[6163]<=16'd4816; ROM2[6163]<=16'd0; ROM3[6163]<=16'd23805; ROM4[6163]<=16'd57294;
ROM1[6164]<=16'd4827; ROM2[6164]<=16'd0; ROM3[6164]<=16'd23789; ROM4[6164]<=16'd57281;
ROM1[6165]<=16'd4849; ROM2[6165]<=16'd0; ROM3[6165]<=16'd23770; ROM4[6165]<=16'd57273;
ROM1[6166]<=16'd4858; ROM2[6166]<=16'd0; ROM3[6166]<=16'd23771; ROM4[6166]<=16'd57277;
ROM1[6167]<=16'd4855; ROM2[6167]<=16'd0; ROM3[6167]<=16'd23790; ROM4[6167]<=16'd57288;
ROM1[6168]<=16'd4853; ROM2[6168]<=16'd0; ROM3[6168]<=16'd23815; ROM4[6168]<=16'd57305;
ROM1[6169]<=16'd4839; ROM2[6169]<=16'd0; ROM3[6169]<=16'd23819; ROM4[6169]<=16'd57299;
ROM1[6170]<=16'd4805; ROM2[6170]<=16'd0; ROM3[6170]<=16'd23803; ROM4[6170]<=16'd57281;
ROM1[6171]<=16'd4794; ROM2[6171]<=16'd0; ROM3[6171]<=16'd23791; ROM4[6171]<=16'd57272;
ROM1[6172]<=16'd4806; ROM2[6172]<=16'd0; ROM3[6172]<=16'd23782; ROM4[6172]<=16'd57267;
ROM1[6173]<=16'd4846; ROM2[6173]<=16'd0; ROM3[6173]<=16'd23784; ROM4[6173]<=16'd57278;
ROM1[6174]<=16'd4888; ROM2[6174]<=16'd0; ROM3[6174]<=16'd23804; ROM4[6174]<=16'd57304;
ROM1[6175]<=16'd4881; ROM2[6175]<=16'd0; ROM3[6175]<=16'd23814; ROM4[6175]<=16'd57310;
ROM1[6176]<=16'd4852; ROM2[6176]<=16'd0; ROM3[6176]<=16'd23811; ROM4[6176]<=16'd57302;
ROM1[6177]<=16'd4828; ROM2[6177]<=16'd0; ROM3[6177]<=16'd23805; ROM4[6177]<=16'd57289;
ROM1[6178]<=16'd4801; ROM2[6178]<=16'd0; ROM3[6178]<=16'd23794; ROM4[6178]<=16'd57276;
ROM1[6179]<=16'd4794; ROM2[6179]<=16'd0; ROM3[6179]<=16'd23794; ROM4[6179]<=16'd57272;
ROM1[6180]<=16'd4811; ROM2[6180]<=16'd0; ROM3[6180]<=16'd23795; ROM4[6180]<=16'd57275;
ROM1[6181]<=16'd4838; ROM2[6181]<=16'd0; ROM3[6181]<=16'd23783; ROM4[6181]<=16'd57276;
ROM1[6182]<=16'd4855; ROM2[6182]<=16'd0; ROM3[6182]<=16'd23761; ROM4[6182]<=16'd57263;
ROM1[6183]<=16'd4852; ROM2[6183]<=16'd0; ROM3[6183]<=16'd23759; ROM4[6183]<=16'd57263;
ROM1[6184]<=16'd4840; ROM2[6184]<=16'd0; ROM3[6184]<=16'd23774; ROM4[6184]<=16'd57270;
ROM1[6185]<=16'd4826; ROM2[6185]<=16'd0; ROM3[6185]<=16'd23790; ROM4[6185]<=16'd57274;
ROM1[6186]<=16'd4815; ROM2[6186]<=16'd0; ROM3[6186]<=16'd23797; ROM4[6186]<=16'd57280;
ROM1[6187]<=16'd4803; ROM2[6187]<=16'd0; ROM3[6187]<=16'd23800; ROM4[6187]<=16'd57281;
ROM1[6188]<=16'd4811; ROM2[6188]<=16'd0; ROM3[6188]<=16'd23797; ROM4[6188]<=16'd57281;
ROM1[6189]<=16'd4832; ROM2[6189]<=16'd0; ROM3[6189]<=16'd23782; ROM4[6189]<=16'd57278;
ROM1[6190]<=16'd4862; ROM2[6190]<=16'd0; ROM3[6190]<=16'd23767; ROM4[6190]<=16'd57276;
ROM1[6191]<=16'd4869; ROM2[6191]<=16'd0; ROM3[6191]<=16'd23763; ROM4[6191]<=16'd57277;
ROM1[6192]<=16'd4850; ROM2[6192]<=16'd0; ROM3[6192]<=16'd23763; ROM4[6192]<=16'd57274;
ROM1[6193]<=16'd4833; ROM2[6193]<=16'd0; ROM3[6193]<=16'd23773; ROM4[6193]<=16'd57273;
ROM1[6194]<=16'd4813; ROM2[6194]<=16'd0; ROM3[6194]<=16'd23773; ROM4[6194]<=16'd57267;
ROM1[6195]<=16'd4797; ROM2[6195]<=16'd0; ROM3[6195]<=16'd23777; ROM4[6195]<=16'd57262;
ROM1[6196]<=16'd4797; ROM2[6196]<=16'd0; ROM3[6196]<=16'd23784; ROM4[6196]<=16'd57265;
ROM1[6197]<=16'd4813; ROM2[6197]<=16'd0; ROM3[6197]<=16'd23780; ROM4[6197]<=16'd57266;
ROM1[6198]<=16'd4856; ROM2[6198]<=16'd0; ROM3[6198]<=16'd23780; ROM4[6198]<=16'd57275;
ROM1[6199]<=16'd4879; ROM2[6199]<=16'd0; ROM3[6199]<=16'd23785; ROM4[6199]<=16'd57285;
ROM1[6200]<=16'd4867; ROM2[6200]<=16'd0; ROM3[6200]<=16'd23788; ROM4[6200]<=16'd57282;
ROM1[6201]<=16'd4834; ROM2[6201]<=16'd0; ROM3[6201]<=16'd23781; ROM4[6201]<=16'd57268;
ROM1[6202]<=16'd4814; ROM2[6202]<=16'd0; ROM3[6202]<=16'd23787; ROM4[6202]<=16'd57266;
ROM1[6203]<=16'd4804; ROM2[6203]<=16'd0; ROM3[6203]<=16'd23798; ROM4[6203]<=16'd57268;
ROM1[6204]<=16'd4801; ROM2[6204]<=16'd0; ROM3[6204]<=16'd23804; ROM4[6204]<=16'd57275;
ROM1[6205]<=16'd4816; ROM2[6205]<=16'd0; ROM3[6205]<=16'd23807; ROM4[6205]<=16'd57280;
ROM1[6206]<=16'd4851; ROM2[6206]<=16'd0; ROM3[6206]<=16'd23797; ROM4[6206]<=16'd57283;
ROM1[6207]<=16'd4878; ROM2[6207]<=16'd0; ROM3[6207]<=16'd23778; ROM4[6207]<=16'd57283;
ROM1[6208]<=16'd4886; ROM2[6208]<=16'd0; ROM3[6208]<=16'd23784; ROM4[6208]<=16'd57290;
ROM1[6209]<=16'd4874; ROM2[6209]<=16'd0; ROM3[6209]<=16'd23795; ROM4[6209]<=16'd57296;
ROM1[6210]<=16'd4834; ROM2[6210]<=16'd0; ROM3[6210]<=16'd23785; ROM4[6210]<=16'd57280;
ROM1[6211]<=16'd4810; ROM2[6211]<=16'd0; ROM3[6211]<=16'd23782; ROM4[6211]<=16'd57269;
ROM1[6212]<=16'd4800; ROM2[6212]<=16'd0; ROM3[6212]<=16'd23787; ROM4[6212]<=16'd57273;
ROM1[6213]<=16'd4820; ROM2[6213]<=16'd0; ROM3[6213]<=16'd23799; ROM4[6213]<=16'd57287;
ROM1[6214]<=16'd4858; ROM2[6214]<=16'd0; ROM3[6214]<=16'd23804; ROM4[6214]<=16'd57298;
ROM1[6215]<=16'd4884; ROM2[6215]<=16'd0; ROM3[6215]<=16'd23786; ROM4[6215]<=16'd57293;
ROM1[6216]<=16'd4887; ROM2[6216]<=16'd0; ROM3[6216]<=16'd23784; ROM4[6216]<=16'd57292;
ROM1[6217]<=16'd4865; ROM2[6217]<=16'd0; ROM3[6217]<=16'd23788; ROM4[6217]<=16'd57290;
ROM1[6218]<=16'd4837; ROM2[6218]<=16'd0; ROM3[6218]<=16'd23790; ROM4[6218]<=16'd57283;
ROM1[6219]<=16'd4829; ROM2[6219]<=16'd0; ROM3[6219]<=16'd23804; ROM4[6219]<=16'd57290;
ROM1[6220]<=16'd4821; ROM2[6220]<=16'd0; ROM3[6220]<=16'd23809; ROM4[6220]<=16'd57291;
ROM1[6221]<=16'd4818; ROM2[6221]<=16'd0; ROM3[6221]<=16'd23801; ROM4[6221]<=16'd57284;
ROM1[6222]<=16'd4823; ROM2[6222]<=16'd0; ROM3[6222]<=16'd23780; ROM4[6222]<=16'd57273;
ROM1[6223]<=16'd4859; ROM2[6223]<=16'd0; ROM3[6223]<=16'd23769; ROM4[6223]<=16'd57276;
ROM1[6224]<=16'd4862; ROM2[6224]<=16'd0; ROM3[6224]<=16'd23750; ROM4[6224]<=16'd57262;
ROM1[6225]<=16'd4826; ROM2[6225]<=16'd0; ROM3[6225]<=16'd23727; ROM4[6225]<=16'd57235;
ROM1[6226]<=16'd4818; ROM2[6226]<=16'd0; ROM3[6226]<=16'd23743; ROM4[6226]<=16'd57245;
ROM1[6227]<=16'd4808; ROM2[6227]<=16'd0; ROM3[6227]<=16'd23753; ROM4[6227]<=16'd57249;
ROM1[6228]<=16'd4792; ROM2[6228]<=16'd0; ROM3[6228]<=16'd23757; ROM4[6228]<=16'd57251;
ROM1[6229]<=16'd4795; ROM2[6229]<=16'd0; ROM3[6229]<=16'd23769; ROM4[6229]<=16'd57258;
ROM1[6230]<=16'd4807; ROM2[6230]<=16'd0; ROM3[6230]<=16'd23768; ROM4[6230]<=16'd57255;
ROM1[6231]<=16'd4829; ROM2[6231]<=16'd0; ROM3[6231]<=16'd23753; ROM4[6231]<=16'd57250;
ROM1[6232]<=16'd4844; ROM2[6232]<=16'd0; ROM3[6232]<=16'd23734; ROM4[6232]<=16'd57242;
ROM1[6233]<=16'd4846; ROM2[6233]<=16'd0; ROM3[6233]<=16'd23740; ROM4[6233]<=16'd57253;
ROM1[6234]<=16'd4852; ROM2[6234]<=16'd0; ROM3[6234]<=16'd23763; ROM4[6234]<=16'd57273;
ROM1[6235]<=16'd4837; ROM2[6235]<=16'd0; ROM3[6235]<=16'd23772; ROM4[6235]<=16'd57274;
ROM1[6236]<=16'd4819; ROM2[6236]<=16'd0; ROM3[6236]<=16'd23771; ROM4[6236]<=16'd57271;
ROM1[6237]<=16'd4820; ROM2[6237]<=16'd0; ROM3[6237]<=16'd23789; ROM4[6237]<=16'd57283;
ROM1[6238]<=16'd4822; ROM2[6238]<=16'd0; ROM3[6238]<=16'd23789; ROM4[6238]<=16'd57282;
ROM1[6239]<=16'd4819; ROM2[6239]<=16'd0; ROM3[6239]<=16'd23757; ROM4[6239]<=16'd57257;
ROM1[6240]<=16'd4838; ROM2[6240]<=16'd0; ROM3[6240]<=16'd23735; ROM4[6240]<=16'd57244;
ROM1[6241]<=16'd4840; ROM2[6241]<=16'd0; ROM3[6241]<=16'd23730; ROM4[6241]<=16'd57239;
ROM1[6242]<=16'd4816; ROM2[6242]<=16'd0; ROM3[6242]<=16'd23731; ROM4[6242]<=16'd57233;
ROM1[6243]<=16'd4806; ROM2[6243]<=16'd0; ROM3[6243]<=16'd23751; ROM4[6243]<=16'd57245;
ROM1[6244]<=16'd4802; ROM2[6244]<=16'd0; ROM3[6244]<=16'd23767; ROM4[6244]<=16'd57257;
ROM1[6245]<=16'd4784; ROM2[6245]<=16'd0; ROM3[6245]<=16'd23770; ROM4[6245]<=16'd57253;
ROM1[6246]<=16'd4792; ROM2[6246]<=16'd0; ROM3[6246]<=16'd23781; ROM4[6246]<=16'd57262;
ROM1[6247]<=16'd4820; ROM2[6247]<=16'd0; ROM3[6247]<=16'd23783; ROM4[6247]<=16'd57267;
ROM1[6248]<=16'd4857; ROM2[6248]<=16'd0; ROM3[6248]<=16'd23776; ROM4[6248]<=16'd57267;
ROM1[6249]<=16'd4875; ROM2[6249]<=16'd0; ROM3[6249]<=16'd23773; ROM4[6249]<=16'd57274;
ROM1[6250]<=16'd4847; ROM2[6250]<=16'd0; ROM3[6250]<=16'd23758; ROM4[6250]<=16'd57259;
ROM1[6251]<=16'd4829; ROM2[6251]<=16'd0; ROM3[6251]<=16'd23766; ROM4[6251]<=16'd57257;
ROM1[6252]<=16'd4816; ROM2[6252]<=16'd0; ROM3[6252]<=16'd23775; ROM4[6252]<=16'd57263;
ROM1[6253]<=16'd4802; ROM2[6253]<=16'd0; ROM3[6253]<=16'd23776; ROM4[6253]<=16'd57263;
ROM1[6254]<=16'd4810; ROM2[6254]<=16'd0; ROM3[6254]<=16'd23790; ROM4[6254]<=16'd57277;
ROM1[6255]<=16'd4827; ROM2[6255]<=16'd0; ROM3[6255]<=16'd23791; ROM4[6255]<=16'd57281;
ROM1[6256]<=16'd4852; ROM2[6256]<=16'd0; ROM3[6256]<=16'd23779; ROM4[6256]<=16'd57276;
ROM1[6257]<=16'd4872; ROM2[6257]<=16'd0; ROM3[6257]<=16'd23763; ROM4[6257]<=16'd57277;
ROM1[6258]<=16'd4870; ROM2[6258]<=16'd0; ROM3[6258]<=16'd23766; ROM4[6258]<=16'd57282;
ROM1[6259]<=16'd4850; ROM2[6259]<=16'd0; ROM3[6259]<=16'd23774; ROM4[6259]<=16'd57284;
ROM1[6260]<=16'd4831; ROM2[6260]<=16'd0; ROM3[6260]<=16'd23777; ROM4[6260]<=16'd57281;
ROM1[6261]<=16'd4810; ROM2[6261]<=16'd0; ROM3[6261]<=16'd23771; ROM4[6261]<=16'd57267;
ROM1[6262]<=16'd4800; ROM2[6262]<=16'd0; ROM3[6262]<=16'd23776; ROM4[6262]<=16'd57270;
ROM1[6263]<=16'd4819; ROM2[6263]<=16'd0; ROM3[6263]<=16'd23791; ROM4[6263]<=16'd57286;
ROM1[6264]<=16'd4828; ROM2[6264]<=16'd0; ROM3[6264]<=16'd23771; ROM4[6264]<=16'd57273;
ROM1[6265]<=16'd4841; ROM2[6265]<=16'd0; ROM3[6265]<=16'd23749; ROM4[6265]<=16'd57258;
ROM1[6266]<=16'd4842; ROM2[6266]<=16'd0; ROM3[6266]<=16'd23744; ROM4[6266]<=16'd57255;
ROM1[6267]<=16'd4822; ROM2[6267]<=16'd0; ROM3[6267]<=16'd23746; ROM4[6267]<=16'd57254;
ROM1[6268]<=16'd4816; ROM2[6268]<=16'd0; ROM3[6268]<=16'd23764; ROM4[6268]<=16'd57267;
ROM1[6269]<=16'd4818; ROM2[6269]<=16'd0; ROM3[6269]<=16'd23782; ROM4[6269]<=16'd57278;
ROM1[6270]<=16'd4798; ROM2[6270]<=16'd0; ROM3[6270]<=16'd23781; ROM4[6270]<=16'd57273;
ROM1[6271]<=16'd4782; ROM2[6271]<=16'd0; ROM3[6271]<=16'd23765; ROM4[6271]<=16'd57259;
ROM1[6272]<=16'd4803; ROM2[6272]<=16'd0; ROM3[6272]<=16'd23763; ROM4[6272]<=16'd57262;
ROM1[6273]<=16'd4844; ROM2[6273]<=16'd0; ROM3[6273]<=16'd23763; ROM4[6273]<=16'd57271;
ROM1[6274]<=16'd4862; ROM2[6274]<=16'd0; ROM3[6274]<=16'd23756; ROM4[6274]<=16'd57266;
ROM1[6275]<=16'd4847; ROM2[6275]<=16'd0; ROM3[6275]<=16'd23760; ROM4[6275]<=16'd57262;
ROM1[6276]<=16'd4841; ROM2[6276]<=16'd0; ROM3[6276]<=16'd23780; ROM4[6276]<=16'd57273;
ROM1[6277]<=16'd4841; ROM2[6277]<=16'd0; ROM3[6277]<=16'd23797; ROM4[6277]<=16'd57286;
ROM1[6278]<=16'd4804; ROM2[6278]<=16'd0; ROM3[6278]<=16'd23779; ROM4[6278]<=16'd57267;
ROM1[6279]<=16'd4797; ROM2[6279]<=16'd0; ROM3[6279]<=16'd23779; ROM4[6279]<=16'd57266;
ROM1[6280]<=16'd4817; ROM2[6280]<=16'd0; ROM3[6280]<=16'd23785; ROM4[6280]<=16'd57279;
ROM1[6281]<=16'd4823; ROM2[6281]<=16'd0; ROM3[6281]<=16'd23753; ROM4[6281]<=16'd57258;
ROM1[6282]<=16'd4845; ROM2[6282]<=16'd0; ROM3[6282]<=16'd23737; ROM4[6282]<=16'd57256;
ROM1[6283]<=16'd4852; ROM2[6283]<=16'd0; ROM3[6283]<=16'd23744; ROM4[6283]<=16'd57267;
ROM1[6284]<=16'd4838; ROM2[6284]<=16'd0; ROM3[6284]<=16'd23750; ROM4[6284]<=16'd57268;
ROM1[6285]<=16'd4824; ROM2[6285]<=16'd0; ROM3[6285]<=16'd23760; ROM4[6285]<=16'd57269;
ROM1[6286]<=16'd4822; ROM2[6286]<=16'd0; ROM3[6286]<=16'd23779; ROM4[6286]<=16'd57282;
ROM1[6287]<=16'd4811; ROM2[6287]<=16'd0; ROM3[6287]<=16'd23785; ROM4[6287]<=16'd57286;
ROM1[6288]<=16'd4810; ROM2[6288]<=16'd0; ROM3[6288]<=16'd23785; ROM4[6288]<=16'd57286;
ROM1[6289]<=16'd4847; ROM2[6289]<=16'd0; ROM3[6289]<=16'd23790; ROM4[6289]<=16'd57298;
ROM1[6290]<=16'd4888; ROM2[6290]<=16'd0; ROM3[6290]<=16'd23793; ROM4[6290]<=16'd57307;
ROM1[6291]<=16'd4888; ROM2[6291]<=16'd0; ROM3[6291]<=16'd23791; ROM4[6291]<=16'd57303;
ROM1[6292]<=16'd4861; ROM2[6292]<=16'd0; ROM3[6292]<=16'd23780; ROM4[6292]<=16'd57285;
ROM1[6293]<=16'd4835; ROM2[6293]<=16'd0; ROM3[6293]<=16'd23779; ROM4[6293]<=16'd57276;
ROM1[6294]<=16'd4821; ROM2[6294]<=16'd0; ROM3[6294]<=16'd23789; ROM4[6294]<=16'd57279;
ROM1[6295]<=16'd4805; ROM2[6295]<=16'd0; ROM3[6295]<=16'd23798; ROM4[6295]<=16'd57278;
ROM1[6296]<=16'd4805; ROM2[6296]<=16'd0; ROM3[6296]<=16'd23806; ROM4[6296]<=16'd57287;
ROM1[6297]<=16'd4836; ROM2[6297]<=16'd0; ROM3[6297]<=16'd23817; ROM4[6297]<=16'd57305;
ROM1[6298]<=16'd4894; ROM2[6298]<=16'd0; ROM3[6298]<=16'd23823; ROM4[6298]<=16'd57324;
ROM1[6299]<=16'd4906; ROM2[6299]<=16'd0; ROM3[6299]<=16'd23804; ROM4[6299]<=16'd57317;
ROM1[6300]<=16'd4873; ROM2[6300]<=16'd0; ROM3[6300]<=16'd23791; ROM4[6300]<=16'd57296;
ROM1[6301]<=16'd4858; ROM2[6301]<=16'd0; ROM3[6301]<=16'd23805; ROM4[6301]<=16'd57301;
ROM1[6302]<=16'd4843; ROM2[6302]<=16'd0; ROM3[6302]<=16'd23810; ROM4[6302]<=16'd57299;
ROM1[6303]<=16'd4816; ROM2[6303]<=16'd0; ROM3[6303]<=16'd23806; ROM4[6303]<=16'd57287;
ROM1[6304]<=16'd4805; ROM2[6304]<=16'd0; ROM3[6304]<=16'd23809; ROM4[6304]<=16'd57286;
ROM1[6305]<=16'd4803; ROM2[6305]<=16'd0; ROM3[6305]<=16'd23793; ROM4[6305]<=16'd57271;
ROM1[6306]<=16'd4819; ROM2[6306]<=16'd0; ROM3[6306]<=16'd23773; ROM4[6306]<=16'd57263;
ROM1[6307]<=16'd4859; ROM2[6307]<=16'd0; ROM3[6307]<=16'd23778; ROM4[6307]<=16'd57280;
ROM1[6308]<=16'd4866; ROM2[6308]<=16'd0; ROM3[6308]<=16'd23788; ROM4[6308]<=16'd57291;
ROM1[6309]<=16'd4840; ROM2[6309]<=16'd0; ROM3[6309]<=16'd23790; ROM4[6309]<=16'd57290;
ROM1[6310]<=16'd4831; ROM2[6310]<=16'd0; ROM3[6310]<=16'd23805; ROM4[6310]<=16'd57300;
ROM1[6311]<=16'd4834; ROM2[6311]<=16'd0; ROM3[6311]<=16'd23826; ROM4[6311]<=16'd57314;
ROM1[6312]<=16'd4812; ROM2[6312]<=16'd0; ROM3[6312]<=16'd23815; ROM4[6312]<=16'd57302;
ROM1[6313]<=16'd4794; ROM2[6313]<=16'd0; ROM3[6313]<=16'd23788; ROM4[6313]<=16'd57279;
ROM1[6314]<=16'd4800; ROM2[6314]<=16'd0; ROM3[6314]<=16'd23763; ROM4[6314]<=16'd57255;
ROM1[6315]<=16'd4824; ROM2[6315]<=16'd0; ROM3[6315]<=16'd23743; ROM4[6315]<=16'd57247;
ROM1[6316]<=16'd4835; ROM2[6316]<=16'd0; ROM3[6316]<=16'd23744; ROM4[6316]<=16'd57253;
ROM1[6317]<=16'd4819; ROM2[6317]<=16'd0; ROM3[6317]<=16'd23752; ROM4[6317]<=16'd57259;
ROM1[6318]<=16'd4793; ROM2[6318]<=16'd0; ROM3[6318]<=16'd23761; ROM4[6318]<=16'd57260;
ROM1[6319]<=16'd4789; ROM2[6319]<=16'd0; ROM3[6319]<=16'd23779; ROM4[6319]<=16'd57266;
ROM1[6320]<=16'd4789; ROM2[6320]<=16'd0; ROM3[6320]<=16'd23796; ROM4[6320]<=16'd57278;
ROM1[6321]<=16'd4781; ROM2[6321]<=16'd0; ROM3[6321]<=16'd23791; ROM4[6321]<=16'd57274;
ROM1[6322]<=16'd4791; ROM2[6322]<=16'd0; ROM3[6322]<=16'd23778; ROM4[6322]<=16'd57263;
ROM1[6323]<=16'd4814; ROM2[6323]<=16'd0; ROM3[6323]<=16'd23761; ROM4[6323]<=16'd57258;
ROM1[6324]<=16'd4826; ROM2[6324]<=16'd0; ROM3[6324]<=16'd23753; ROM4[6324]<=16'd57256;
ROM1[6325]<=16'd4823; ROM2[6325]<=16'd0; ROM3[6325]<=16'd23770; ROM4[6325]<=16'd57263;
ROM1[6326]<=16'd4814; ROM2[6326]<=16'd0; ROM3[6326]<=16'd23789; ROM4[6326]<=16'd57275;
ROM1[6327]<=16'd4797; ROM2[6327]<=16'd0; ROM3[6327]<=16'd23791; ROM4[6327]<=16'd57270;
ROM1[6328]<=16'd4790; ROM2[6328]<=16'd0; ROM3[6328]<=16'd23797; ROM4[6328]<=16'd57271;
ROM1[6329]<=16'd4803; ROM2[6329]<=16'd0; ROM3[6329]<=16'd23814; ROM4[6329]<=16'd57287;
ROM1[6330]<=16'd4802; ROM2[6330]<=16'd0; ROM3[6330]<=16'd23798; ROM4[6330]<=16'd57278;
ROM1[6331]<=16'd4817; ROM2[6331]<=16'd0; ROM3[6331]<=16'd23779; ROM4[6331]<=16'd57273;
ROM1[6332]<=16'd4838; ROM2[6332]<=16'd0; ROM3[6332]<=16'd23769; ROM4[6332]<=16'd57270;
ROM1[6333]<=16'd4833; ROM2[6333]<=16'd0; ROM3[6333]<=16'd23768; ROM4[6333]<=16'd57268;
ROM1[6334]<=16'd4828; ROM2[6334]<=16'd0; ROM3[6334]<=16'd23786; ROM4[6334]<=16'd57280;
ROM1[6335]<=16'd4831; ROM2[6335]<=16'd0; ROM3[6335]<=16'd23806; ROM4[6335]<=16'd57296;
ROM1[6336]<=16'd4835; ROM2[6336]<=16'd0; ROM3[6336]<=16'd23828; ROM4[6336]<=16'd57313;
ROM1[6337]<=16'd4812; ROM2[6337]<=16'd0; ROM3[6337]<=16'd23820; ROM4[6337]<=16'd57299;
ROM1[6338]<=16'd4803; ROM2[6338]<=16'd0; ROM3[6338]<=16'd23803; ROM4[6338]<=16'd57284;
ROM1[6339]<=16'd4831; ROM2[6339]<=16'd0; ROM3[6339]<=16'd23795; ROM4[6339]<=16'd57288;
ROM1[6340]<=16'd4860; ROM2[6340]<=16'd0; ROM3[6340]<=16'd23777; ROM4[6340]<=16'd57284;
ROM1[6341]<=16'd4859; ROM2[6341]<=16'd0; ROM3[6341]<=16'd23768; ROM4[6341]<=16'd57280;
ROM1[6342]<=16'd4846; ROM2[6342]<=16'd0; ROM3[6342]<=16'd23776; ROM4[6342]<=16'd57284;
ROM1[6343]<=16'd4826; ROM2[6343]<=16'd0; ROM3[6343]<=16'd23785; ROM4[6343]<=16'd57280;
ROM1[6344]<=16'd4804; ROM2[6344]<=16'd0; ROM3[6344]<=16'd23787; ROM4[6344]<=16'd57269;
ROM1[6345]<=16'd4799; ROM2[6345]<=16'd0; ROM3[6345]<=16'd23800; ROM4[6345]<=16'd57275;
ROM1[6346]<=16'd4817; ROM2[6346]<=16'd0; ROM3[6346]<=16'd23819; ROM4[6346]<=16'd57292;
ROM1[6347]<=16'd4843; ROM2[6347]<=16'd0; ROM3[6347]<=16'd23817; ROM4[6347]<=16'd57301;
ROM1[6348]<=16'd4852; ROM2[6348]<=16'd0; ROM3[6348]<=16'd23783; ROM4[6348]<=16'd57280;
ROM1[6349]<=16'd4860; ROM2[6349]<=16'd0; ROM3[6349]<=16'd23765; ROM4[6349]<=16'd57270;
ROM1[6350]<=16'd4857; ROM2[6350]<=16'd0; ROM3[6350]<=16'd23777; ROM4[6350]<=16'd57276;
ROM1[6351]<=16'd4831; ROM2[6351]<=16'd0; ROM3[6351]<=16'd23778; ROM4[6351]<=16'd57266;
ROM1[6352]<=16'd4817; ROM2[6352]<=16'd0; ROM3[6352]<=16'd23788; ROM4[6352]<=16'd57271;
ROM1[6353]<=16'd4808; ROM2[6353]<=16'd0; ROM3[6353]<=16'd23801; ROM4[6353]<=16'd57281;
ROM1[6354]<=16'd4801; ROM2[6354]<=16'd0; ROM3[6354]<=16'd23800; ROM4[6354]<=16'd57281;
ROM1[6355]<=16'd4807; ROM2[6355]<=16'd0; ROM3[6355]<=16'd23797; ROM4[6355]<=16'd57281;
ROM1[6356]<=16'd4831; ROM2[6356]<=16'd0; ROM3[6356]<=16'd23781; ROM4[6356]<=16'd57277;
ROM1[6357]<=16'd4852; ROM2[6357]<=16'd0; ROM3[6357]<=16'd23764; ROM4[6357]<=16'd57274;
ROM1[6358]<=16'd4835; ROM2[6358]<=16'd0; ROM3[6358]<=16'd23756; ROM4[6358]<=16'd57265;
ROM1[6359]<=16'd4826; ROM2[6359]<=16'd0; ROM3[6359]<=16'd23767; ROM4[6359]<=16'd57271;
ROM1[6360]<=16'd4837; ROM2[6360]<=16'd0; ROM3[6360]<=16'd23802; ROM4[6360]<=16'd57299;
ROM1[6361]<=16'd4827; ROM2[6361]<=16'd0; ROM3[6361]<=16'd23808; ROM4[6361]<=16'd57298;
ROM1[6362]<=16'd4814; ROM2[6362]<=16'd0; ROM3[6362]<=16'd23810; ROM4[6362]<=16'd57296;
ROM1[6363]<=16'd4806; ROM2[6363]<=16'd0; ROM3[6363]<=16'd23801; ROM4[6363]<=16'd57288;
ROM1[6364]<=16'd4814; ROM2[6364]<=16'd0; ROM3[6364]<=16'd23782; ROM4[6364]<=16'd57275;
ROM1[6365]<=16'd4850; ROM2[6365]<=16'd0; ROM3[6365]<=16'd23781; ROM4[6365]<=16'd57282;
ROM1[6366]<=16'd4855; ROM2[6366]<=16'd0; ROM3[6366]<=16'd23779; ROM4[6366]<=16'd57284;
ROM1[6367]<=16'd4844; ROM2[6367]<=16'd0; ROM3[6367]<=16'd23789; ROM4[6367]<=16'd57290;
ROM1[6368]<=16'd4834; ROM2[6368]<=16'd0; ROM3[6368]<=16'd23804; ROM4[6368]<=16'd57296;
ROM1[6369]<=16'd4822; ROM2[6369]<=16'd0; ROM3[6369]<=16'd23810; ROM4[6369]<=16'd57297;
ROM1[6370]<=16'd4807; ROM2[6370]<=16'd0; ROM3[6370]<=16'd23809; ROM4[6370]<=16'd57298;
ROM1[6371]<=16'd4805; ROM2[6371]<=16'd0; ROM3[6371]<=16'd23803; ROM4[6371]<=16'd57294;
ROM1[6372]<=16'd4820; ROM2[6372]<=16'd0; ROM3[6372]<=16'd23789; ROM4[6372]<=16'd57288;
ROM1[6373]<=16'd4848; ROM2[6373]<=16'd0; ROM3[6373]<=16'd23772; ROM4[6373]<=16'd57289;
ROM1[6374]<=16'd4874; ROM2[6374]<=16'd0; ROM3[6374]<=16'd23777; ROM4[6374]<=16'd57298;
ROM1[6375]<=16'd4879; ROM2[6375]<=16'd0; ROM3[6375]<=16'd23800; ROM4[6375]<=16'd57314;
ROM1[6376]<=16'd4880; ROM2[6376]<=16'd0; ROM3[6376]<=16'd23827; ROM4[6376]<=16'd57336;
ROM1[6377]<=16'd4866; ROM2[6377]<=16'd0; ROM3[6377]<=16'd23835; ROM4[6377]<=16'd57334;
ROM1[6378]<=16'd4822; ROM2[6378]<=16'd0; ROM3[6378]<=16'd23817; ROM4[6378]<=16'd57307;
ROM1[6379]<=16'd4797; ROM2[6379]<=16'd0; ROM3[6379]<=16'd23804; ROM4[6379]<=16'd57292;
ROM1[6380]<=16'd4801; ROM2[6380]<=16'd0; ROM3[6380]<=16'd23800; ROM4[6380]<=16'd57290;
ROM1[6381]<=16'd4833; ROM2[6381]<=16'd0; ROM3[6381]<=16'd23797; ROM4[6381]<=16'd57295;
ROM1[6382]<=16'd4873; ROM2[6382]<=16'd0; ROM3[6382]<=16'd23802; ROM4[6382]<=16'd57303;
ROM1[6383]<=16'd4866; ROM2[6383]<=16'd0; ROM3[6383]<=16'd23796; ROM4[6383]<=16'd57296;
ROM1[6384]<=16'd4839; ROM2[6384]<=16'd0; ROM3[6384]<=16'd23793; ROM4[6384]<=16'd57287;
ROM1[6385]<=16'd4829; ROM2[6385]<=16'd0; ROM3[6385]<=16'd23811; ROM4[6385]<=16'd57295;
ROM1[6386]<=16'd4828; ROM2[6386]<=16'd0; ROM3[6386]<=16'd23827; ROM4[6386]<=16'd57310;
ROM1[6387]<=16'd4809; ROM2[6387]<=16'd0; ROM3[6387]<=16'd23827; ROM4[6387]<=16'd57305;
ROM1[6388]<=16'd4814; ROM2[6388]<=16'd0; ROM3[6388]<=16'd23830; ROM4[6388]<=16'd57305;
ROM1[6389]<=16'd4836; ROM2[6389]<=16'd0; ROM3[6389]<=16'd23821; ROM4[6389]<=16'd57304;
ROM1[6390]<=16'd4847; ROM2[6390]<=16'd0; ROM3[6390]<=16'd23793; ROM4[6390]<=16'd57287;
ROM1[6391]<=16'd4853; ROM2[6391]<=16'd0; ROM3[6391]<=16'd23791; ROM4[6391]<=16'd57288;
ROM1[6392]<=16'd4832; ROM2[6392]<=16'd0; ROM3[6392]<=16'd23789; ROM4[6392]<=16'd57280;
ROM1[6393]<=16'd4803; ROM2[6393]<=16'd0; ROM3[6393]<=16'd23785; ROM4[6393]<=16'd57270;
ROM1[6394]<=16'd4792; ROM2[6394]<=16'd0; ROM3[6394]<=16'd23791; ROM4[6394]<=16'd57275;
ROM1[6395]<=16'd4773; ROM2[6395]<=16'd0; ROM3[6395]<=16'd23793; ROM4[6395]<=16'd57267;
ROM1[6396]<=16'd4763; ROM2[6396]<=16'd0; ROM3[6396]<=16'd23791; ROM4[6396]<=16'd57263;
ROM1[6397]<=16'd4783; ROM2[6397]<=16'd0; ROM3[6397]<=16'd23784; ROM4[6397]<=16'd57262;
ROM1[6398]<=16'd4822; ROM2[6398]<=16'd0; ROM3[6398]<=16'd23777; ROM4[6398]<=16'd57266;
ROM1[6399]<=16'd4846; ROM2[6399]<=16'd0; ROM3[6399]<=16'd23776; ROM4[6399]<=16'd57280;
ROM1[6400]<=16'd4851; ROM2[6400]<=16'd0; ROM3[6400]<=16'd23792; ROM4[6400]<=16'd57294;
ROM1[6401]<=16'd4834; ROM2[6401]<=16'd0; ROM3[6401]<=16'd23806; ROM4[6401]<=16'd57301;
ROM1[6402]<=16'd4803; ROM2[6402]<=16'd0; ROM3[6402]<=16'd23800; ROM4[6402]<=16'd57288;
ROM1[6403]<=16'd4787; ROM2[6403]<=16'd0; ROM3[6403]<=16'd23809; ROM4[6403]<=16'd57284;
ROM1[6404]<=16'd4778; ROM2[6404]<=16'd0; ROM3[6404]<=16'd23809; ROM4[6404]<=16'd57284;
ROM1[6405]<=16'd4784; ROM2[6405]<=16'd0; ROM3[6405]<=16'd23794; ROM4[6405]<=16'd57275;
ROM1[6406]<=16'd4798; ROM2[6406]<=16'd0; ROM3[6406]<=16'd23771; ROM4[6406]<=16'd57261;
ROM1[6407]<=16'd4816; ROM2[6407]<=16'd0; ROM3[6407]<=16'd23751; ROM4[6407]<=16'd57256;
ROM1[6408]<=16'd4807; ROM2[6408]<=16'd0; ROM3[6408]<=16'd23746; ROM4[6408]<=16'd57252;
ROM1[6409]<=16'd4792; ROM2[6409]<=16'd0; ROM3[6409]<=16'd23754; ROM4[6409]<=16'd57254;
ROM1[6410]<=16'd4784; ROM2[6410]<=16'd0; ROM3[6410]<=16'd23765; ROM4[6410]<=16'd57256;
ROM1[6411]<=16'd4759; ROM2[6411]<=16'd0; ROM3[6411]<=16'd23760; ROM4[6411]<=16'd57245;
ROM1[6412]<=16'd4747; ROM2[6412]<=16'd0; ROM3[6412]<=16'd23763; ROM4[6412]<=16'd57246;
ROM1[6413]<=16'd4762; ROM2[6413]<=16'd0; ROM3[6413]<=16'd23764; ROM4[6413]<=16'd57250;
ROM1[6414]<=16'd4782; ROM2[6414]<=16'd0; ROM3[6414]<=16'd23750; ROM4[6414]<=16'd57246;
ROM1[6415]<=16'd4808; ROM2[6415]<=16'd0; ROM3[6415]<=16'd23732; ROM4[6415]<=16'd57242;
ROM1[6416]<=16'd4807; ROM2[6416]<=16'd0; ROM3[6416]<=16'd23725; ROM4[6416]<=16'd57239;
ROM1[6417]<=16'd4793; ROM2[6417]<=16'd0; ROM3[6417]<=16'd23735; ROM4[6417]<=16'd57241;
ROM1[6418]<=16'd4801; ROM2[6418]<=16'd0; ROM3[6418]<=16'd23766; ROM4[6418]<=16'd57265;
ROM1[6419]<=16'd4804; ROM2[6419]<=16'd0; ROM3[6419]<=16'd23790; ROM4[6419]<=16'd57278;
ROM1[6420]<=16'd4783; ROM2[6420]<=16'd0; ROM3[6420]<=16'd23784; ROM4[6420]<=16'd57272;
ROM1[6421]<=16'd4772; ROM2[6421]<=16'd0; ROM3[6421]<=16'd23773; ROM4[6421]<=16'd57265;
ROM1[6422]<=16'd4784; ROM2[6422]<=16'd0; ROM3[6422]<=16'd23766; ROM4[6422]<=16'd57261;
ROM1[6423]<=16'd4822; ROM2[6423]<=16'd0; ROM3[6423]<=16'd23753; ROM4[6423]<=16'd57266;
ROM1[6424]<=16'd4841; ROM2[6424]<=16'd0; ROM3[6424]<=16'd23745; ROM4[6424]<=16'd57263;
ROM1[6425]<=16'd4831; ROM2[6425]<=16'd0; ROM3[6425]<=16'd23750; ROM4[6425]<=16'd57263;
ROM1[6426]<=16'd4809; ROM2[6426]<=16'd0; ROM3[6426]<=16'd23759; ROM4[6426]<=16'd57266;
ROM1[6427]<=16'd4784; ROM2[6427]<=16'd0; ROM3[6427]<=16'd23768; ROM4[6427]<=16'd57263;
ROM1[6428]<=16'd4783; ROM2[6428]<=16'd0; ROM3[6428]<=16'd23791; ROM4[6428]<=16'd57282;
ROM1[6429]<=16'd4772; ROM2[6429]<=16'd0; ROM3[6429]<=16'd23791; ROM4[6429]<=16'd57278;
ROM1[6430]<=16'd4762; ROM2[6430]<=16'd0; ROM3[6430]<=16'd23763; ROM4[6430]<=16'd57252;
ROM1[6431]<=16'd4795; ROM2[6431]<=16'd0; ROM3[6431]<=16'd23750; ROM4[6431]<=16'd57250;
ROM1[6432]<=16'd4819; ROM2[6432]<=16'd0; ROM3[6432]<=16'd23737; ROM4[6432]<=16'd57247;
ROM1[6433]<=16'd4809; ROM2[6433]<=16'd0; ROM3[6433]<=16'd23733; ROM4[6433]<=16'd57245;
ROM1[6434]<=16'd4802; ROM2[6434]<=16'd0; ROM3[6434]<=16'd23750; ROM4[6434]<=16'd57260;
ROM1[6435]<=16'd4789; ROM2[6435]<=16'd0; ROM3[6435]<=16'd23763; ROM4[6435]<=16'd57268;
ROM1[6436]<=16'd4774; ROM2[6436]<=16'd0; ROM3[6436]<=16'd23766; ROM4[6436]<=16'd57261;
ROM1[6437]<=16'd4760; ROM2[6437]<=16'd0; ROM3[6437]<=16'd23772; ROM4[6437]<=16'd57260;
ROM1[6438]<=16'd4766; ROM2[6438]<=16'd0; ROM3[6438]<=16'd23771; ROM4[6438]<=16'd57262;
ROM1[6439]<=16'd4791; ROM2[6439]<=16'd0; ROM3[6439]<=16'd23762; ROM4[6439]<=16'd57263;
ROM1[6440]<=16'd4815; ROM2[6440]<=16'd0; ROM3[6440]<=16'd23749; ROM4[6440]<=16'd57259;
ROM1[6441]<=16'd4813; ROM2[6441]<=16'd0; ROM3[6441]<=16'd23743; ROM4[6441]<=16'd57258;
ROM1[6442]<=16'd4802; ROM2[6442]<=16'd0; ROM3[6442]<=16'd23756; ROM4[6442]<=16'd57264;
ROM1[6443]<=16'd4785; ROM2[6443]<=16'd0; ROM3[6443]<=16'd23771; ROM4[6443]<=16'd57267;
ROM1[6444]<=16'd4794; ROM2[6444]<=16'd0; ROM3[6444]<=16'd23795; ROM4[6444]<=16'd57290;
ROM1[6445]<=16'd4790; ROM2[6445]<=16'd0; ROM3[6445]<=16'd23805; ROM4[6445]<=16'd57296;
ROM1[6446]<=16'd4767; ROM2[6446]<=16'd0; ROM3[6446]<=16'd23788; ROM4[6446]<=16'd57275;
ROM1[6447]<=16'd4762; ROM2[6447]<=16'd0; ROM3[6447]<=16'd23764; ROM4[6447]<=16'd57256;
ROM1[6448]<=16'd4777; ROM2[6448]<=16'd0; ROM3[6448]<=16'd23740; ROM4[6448]<=16'd57243;
ROM1[6449]<=16'd4812; ROM2[6449]<=16'd0; ROM3[6449]<=16'd23750; ROM4[6449]<=16'd57260;
ROM1[6450]<=16'd4814; ROM2[6450]<=16'd0; ROM3[6450]<=16'd23761; ROM4[6450]<=16'd57268;
ROM1[6451]<=16'd4796; ROM2[6451]<=16'd0; ROM3[6451]<=16'd23763; ROM4[6451]<=16'd57265;
ROM1[6452]<=16'd4786; ROM2[6452]<=16'd0; ROM3[6452]<=16'd23771; ROM4[6452]<=16'd57268;
ROM1[6453]<=16'd4782; ROM2[6453]<=16'd0; ROM3[6453]<=16'd23792; ROM4[6453]<=16'd57280;
ROM1[6454]<=16'd4778; ROM2[6454]<=16'd0; ROM3[6454]<=16'd23796; ROM4[6454]<=16'd57284;
ROM1[6455]<=16'd4783; ROM2[6455]<=16'd0; ROM3[6455]<=16'd23786; ROM4[6455]<=16'd57278;
ROM1[6456]<=16'd4819; ROM2[6456]<=16'd0; ROM3[6456]<=16'd23787; ROM4[6456]<=16'd57285;
ROM1[6457]<=16'd4847; ROM2[6457]<=16'd0; ROM3[6457]<=16'd23775; ROM4[6457]<=16'd57285;
ROM1[6458]<=16'd4832; ROM2[6458]<=16'd0; ROM3[6458]<=16'd23766; ROM4[6458]<=16'd57276;
ROM1[6459]<=16'd4818; ROM2[6459]<=16'd0; ROM3[6459]<=16'd23775; ROM4[6459]<=16'd57278;
ROM1[6460]<=16'd4803; ROM2[6460]<=16'd0; ROM3[6460]<=16'd23782; ROM4[6460]<=16'd57280;
ROM1[6461]<=16'd4772; ROM2[6461]<=16'd0; ROM3[6461]<=16'd23773; ROM4[6461]<=16'd57265;
ROM1[6462]<=16'd4760; ROM2[6462]<=16'd0; ROM3[6462]<=16'd23772; ROM4[6462]<=16'd57263;
ROM1[6463]<=16'd4773; ROM2[6463]<=16'd0; ROM3[6463]<=16'd23771; ROM4[6463]<=16'd57264;
ROM1[6464]<=16'd4787; ROM2[6464]<=16'd0; ROM3[6464]<=16'd23751; ROM4[6464]<=16'd57249;
ROM1[6465]<=16'd4808; ROM2[6465]<=16'd0; ROM3[6465]<=16'd23733; ROM4[6465]<=16'd57242;
ROM1[6466]<=16'd4820; ROM2[6466]<=16'd0; ROM3[6466]<=16'd23744; ROM4[6466]<=16'd57255;
ROM1[6467]<=16'd4817; ROM2[6467]<=16'd0; ROM3[6467]<=16'd23765; ROM4[6467]<=16'd57273;
ROM1[6468]<=16'd4804; ROM2[6468]<=16'd0; ROM3[6468]<=16'd23773; ROM4[6468]<=16'd57277;
ROM1[6469]<=16'd4785; ROM2[6469]<=16'd0; ROM3[6469]<=16'd23771; ROM4[6469]<=16'd57269;
ROM1[6470]<=16'd4766; ROM2[6470]<=16'd0; ROM3[6470]<=16'd23773; ROM4[6470]<=16'd57267;
ROM1[6471]<=16'd4764; ROM2[6471]<=16'd0; ROM3[6471]<=16'd23775; ROM4[6471]<=16'd57269;
ROM1[6472]<=16'd4774; ROM2[6472]<=16'd0; ROM3[6472]<=16'd23765; ROM4[6472]<=16'd57265;
ROM1[6473]<=16'd4813; ROM2[6473]<=16'd0; ROM3[6473]<=16'd23760; ROM4[6473]<=16'd57270;
ROM1[6474]<=16'd4841; ROM2[6474]<=16'd0; ROM3[6474]<=16'd23761; ROM4[6474]<=16'd57276;
ROM1[6475]<=16'd4824; ROM2[6475]<=16'd0; ROM3[6475]<=16'd23755; ROM4[6475]<=16'd57270;
ROM1[6476]<=16'd4799; ROM2[6476]<=16'd0; ROM3[6476]<=16'd23758; ROM4[6476]<=16'd57264;
ROM1[6477]<=16'd4797; ROM2[6477]<=16'd0; ROM3[6477]<=16'd23772; ROM4[6477]<=16'd57274;
ROM1[6478]<=16'd4799; ROM2[6478]<=16'd0; ROM3[6478]<=16'd23785; ROM4[6478]<=16'd57286;
ROM1[6479]<=16'd4788; ROM2[6479]<=16'd0; ROM3[6479]<=16'd23786; ROM4[6479]<=16'd57279;
ROM1[6480]<=16'd4790; ROM2[6480]<=16'd0; ROM3[6480]<=16'd23775; ROM4[6480]<=16'd57273;
ROM1[6481]<=16'd4822; ROM2[6481]<=16'd0; ROM3[6481]<=16'd23768; ROM4[6481]<=16'd57277;
ROM1[6482]<=16'd4852; ROM2[6482]<=16'd0; ROM3[6482]<=16'd23765; ROM4[6482]<=16'd57281;
ROM1[6483]<=16'd4850; ROM2[6483]<=16'd0; ROM3[6483]<=16'd23769; ROM4[6483]<=16'd57285;
ROM1[6484]<=16'd4818; ROM2[6484]<=16'd0; ROM3[6484]<=16'd23758; ROM4[6484]<=16'd57271;
ROM1[6485]<=16'd4787; ROM2[6485]<=16'd0; ROM3[6485]<=16'd23747; ROM4[6485]<=16'd57256;
ROM1[6486]<=16'd4765; ROM2[6486]<=16'd0; ROM3[6486]<=16'd23743; ROM4[6486]<=16'd57246;
ROM1[6487]<=16'd4752; ROM2[6487]<=16'd0; ROM3[6487]<=16'd23750; ROM4[6487]<=16'd57247;
ROM1[6488]<=16'd4776; ROM2[6488]<=16'd0; ROM3[6488]<=16'd23769; ROM4[6488]<=16'd57266;
ROM1[6489]<=16'd4808; ROM2[6489]<=16'd0; ROM3[6489]<=16'd23772; ROM4[6489]<=16'd57271;
ROM1[6490]<=16'd4825; ROM2[6490]<=16'd0; ROM3[6490]<=16'd23755; ROM4[6490]<=16'd57266;
ROM1[6491]<=16'd4827; ROM2[6491]<=16'd0; ROM3[6491]<=16'd23755; ROM4[6491]<=16'd57273;
ROM1[6492]<=16'd4811; ROM2[6492]<=16'd0; ROM3[6492]<=16'd23765; ROM4[6492]<=16'd57272;
ROM1[6493]<=16'd4796; ROM2[6493]<=16'd0; ROM3[6493]<=16'd23782; ROM4[6493]<=16'd57283;
ROM1[6494]<=16'd4783; ROM2[6494]<=16'd0; ROM3[6494]<=16'd23785; ROM4[6494]<=16'd57285;
ROM1[6495]<=16'd4761; ROM2[6495]<=16'd0; ROM3[6495]<=16'd23773; ROM4[6495]<=16'd57268;
ROM1[6496]<=16'd4750; ROM2[6496]<=16'd0; ROM3[6496]<=16'd23763; ROM4[6496]<=16'd57259;
ROM1[6497]<=16'd4756; ROM2[6497]<=16'd0; ROM3[6497]<=16'd23745; ROM4[6497]<=16'd57251;
ROM1[6498]<=16'd4793; ROM2[6498]<=16'd0; ROM3[6498]<=16'd23739; ROM4[6498]<=16'd57256;
ROM1[6499]<=16'd4821; ROM2[6499]<=16'd0; ROM3[6499]<=16'd23747; ROM4[6499]<=16'd57269;
ROM1[6500]<=16'd4812; ROM2[6500]<=16'd0; ROM3[6500]<=16'd23754; ROM4[6500]<=16'd57271;
ROM1[6501]<=16'd4794; ROM2[6501]<=16'd0; ROM3[6501]<=16'd23762; ROM4[6501]<=16'd57271;
ROM1[6502]<=16'd4798; ROM2[6502]<=16'd0; ROM3[6502]<=16'd23791; ROM4[6502]<=16'd57292;
ROM1[6503]<=16'd4787; ROM2[6503]<=16'd0; ROM3[6503]<=16'd23801; ROM4[6503]<=16'd57296;
ROM1[6504]<=16'd4760; ROM2[6504]<=16'd0; ROM3[6504]<=16'd23778; ROM4[6504]<=16'd57273;
ROM1[6505]<=16'd4762; ROM2[6505]<=16'd0; ROM3[6505]<=16'd23761; ROM4[6505]<=16'd57258;
ROM1[6506]<=16'd4788; ROM2[6506]<=16'd0; ROM3[6506]<=16'd23742; ROM4[6506]<=16'd57250;
ROM1[6507]<=16'd4810; ROM2[6507]<=16'd0; ROM3[6507]<=16'd23728; ROM4[6507]<=16'd57246;
ROM1[6508]<=16'd4811; ROM2[6508]<=16'd0; ROM3[6508]<=16'd23742; ROM4[6508]<=16'd57257;
ROM1[6509]<=16'd4797; ROM2[6509]<=16'd0; ROM3[6509]<=16'd23759; ROM4[6509]<=16'd57265;
ROM1[6510]<=16'd4767; ROM2[6510]<=16'd0; ROM3[6510]<=16'd23757; ROM4[6510]<=16'd57252;
ROM1[6511]<=16'd4749; ROM2[6511]<=16'd0; ROM3[6511]<=16'd23758; ROM4[6511]<=16'd57245;
ROM1[6512]<=16'd4748; ROM2[6512]<=16'd0; ROM3[6512]<=16'd23770; ROM4[6512]<=16'd57254;
ROM1[6513]<=16'd4752; ROM2[6513]<=16'd0; ROM3[6513]<=16'd23771; ROM4[6513]<=16'd57257;
ROM1[6514]<=16'd4775; ROM2[6514]<=16'd0; ROM3[6514]<=16'd23767; ROM4[6514]<=16'd57260;
ROM1[6515]<=16'd4808; ROM2[6515]<=16'd0; ROM3[6515]<=16'd23757; ROM4[6515]<=16'd57265;
ROM1[6516]<=16'd4818; ROM2[6516]<=16'd0; ROM3[6516]<=16'd23758; ROM4[6516]<=16'd57268;
ROM1[6517]<=16'd4812; ROM2[6517]<=16'd0; ROM3[6517]<=16'd23768; ROM4[6517]<=16'd57274;
ROM1[6518]<=16'd4799; ROM2[6518]<=16'd0; ROM3[6518]<=16'd23779; ROM4[6518]<=16'd57277;
ROM1[6519]<=16'd4783; ROM2[6519]<=16'd0; ROM3[6519]<=16'd23783; ROM4[6519]<=16'd57276;
ROM1[6520]<=16'd4767; ROM2[6520]<=16'd0; ROM3[6520]<=16'd23786; ROM4[6520]<=16'd57272;
ROM1[6521]<=16'd4766; ROM2[6521]<=16'd0; ROM3[6521]<=16'd23781; ROM4[6521]<=16'd57268;
ROM1[6522]<=16'd4778; ROM2[6522]<=16'd0; ROM3[6522]<=16'd23769; ROM4[6522]<=16'd57266;
ROM1[6523]<=16'd4817; ROM2[6523]<=16'd0; ROM3[6523]<=16'd23770; ROM4[6523]<=16'd57276;
ROM1[6524]<=16'd4843; ROM2[6524]<=16'd0; ROM3[6524]<=16'd23778; ROM4[6524]<=16'd57290;
ROM1[6525]<=16'd4835; ROM2[6525]<=16'd0; ROM3[6525]<=16'd23792; ROM4[6525]<=16'd57301;
ROM1[6526]<=16'd4808; ROM2[6526]<=16'd0; ROM3[6526]<=16'd23794; ROM4[6526]<=16'd57296;
ROM1[6527]<=16'd4780; ROM2[6527]<=16'd0; ROM3[6527]<=16'd23786; ROM4[6527]<=16'd57278;
ROM1[6528]<=16'd4772; ROM2[6528]<=16'd0; ROM3[6528]<=16'd23801; ROM4[6528]<=16'd57288;
ROM1[6529]<=16'd4763; ROM2[6529]<=16'd0; ROM3[6529]<=16'd23804; ROM4[6529]<=16'd57288;
ROM1[6530]<=16'd4777; ROM2[6530]<=16'd0; ROM3[6530]<=16'd23804; ROM4[6530]<=16'd57285;
ROM1[6531]<=16'd4818; ROM2[6531]<=16'd0; ROM3[6531]<=16'd23804; ROM4[6531]<=16'd57297;
ROM1[6532]<=16'd4835; ROM2[6532]<=16'd0; ROM3[6532]<=16'd23787; ROM4[6532]<=16'd57288;
ROM1[6533]<=16'd4828; ROM2[6533]<=16'd0; ROM3[6533]<=16'd23787; ROM4[6533]<=16'd57284;
ROM1[6534]<=16'd4826; ROM2[6534]<=16'd0; ROM3[6534]<=16'd23806; ROM4[6534]<=16'd57297;
ROM1[6535]<=16'd4810; ROM2[6535]<=16'd0; ROM3[6535]<=16'd23817; ROM4[6535]<=16'd57300;
ROM1[6536]<=16'd4781; ROM2[6536]<=16'd0; ROM3[6536]<=16'd23805; ROM4[6536]<=16'd57289;
ROM1[6537]<=16'd4763; ROM2[6537]<=16'd0; ROM3[6537]<=16'd23802; ROM4[6537]<=16'd57284;
ROM1[6538]<=16'd4764; ROM2[6538]<=16'd0; ROM3[6538]<=16'd23798; ROM4[6538]<=16'd57282;
ROM1[6539]<=16'd4776; ROM2[6539]<=16'd0; ROM3[6539]<=16'd23773; ROM4[6539]<=16'd57267;
ROM1[6540]<=16'd4810; ROM2[6540]<=16'd0; ROM3[6540]<=16'd23766; ROM4[6540]<=16'd57270;
ROM1[6541]<=16'd4832; ROM2[6541]<=16'd0; ROM3[6541]<=16'd23778; ROM4[6541]<=16'd57284;
ROM1[6542]<=16'd4822; ROM2[6542]<=16'd0; ROM3[6542]<=16'd23788; ROM4[6542]<=16'd57292;
ROM1[6543]<=16'd4796; ROM2[6543]<=16'd0; ROM3[6543]<=16'd23790; ROM4[6543]<=16'd57287;
ROM1[6544]<=16'd4769; ROM2[6544]<=16'd0; ROM3[6544]<=16'd23782; ROM4[6544]<=16'd57272;
ROM1[6545]<=16'd4741; ROM2[6545]<=16'd0; ROM3[6545]<=16'd23774; ROM4[6545]<=16'd57259;
ROM1[6546]<=16'd4730; ROM2[6546]<=16'd0; ROM3[6546]<=16'd23763; ROM4[6546]<=16'd57249;
ROM1[6547]<=16'd4756; ROM2[6547]<=16'd0; ROM3[6547]<=16'd23771; ROM4[6547]<=16'd57256;
ROM1[6548]<=16'd4816; ROM2[6548]<=16'd0; ROM3[6548]<=16'd23787; ROM4[6548]<=16'd57284;
ROM1[6549]<=16'd4833; ROM2[6549]<=16'd0; ROM3[6549]<=16'd23783; ROM4[6549]<=16'd57289;
ROM1[6550]<=16'd4796; ROM2[6550]<=16'd0; ROM3[6550]<=16'd23768; ROM4[6550]<=16'd57270;
ROM1[6551]<=16'd4769; ROM2[6551]<=16'd0; ROM3[6551]<=16'd23771; ROM4[6551]<=16'd57266;
ROM1[6552]<=16'd4747; ROM2[6552]<=16'd0; ROM3[6552]<=16'd23770; ROM4[6552]<=16'd57258;
ROM1[6553]<=16'd4732; ROM2[6553]<=16'd0; ROM3[6553]<=16'd23776; ROM4[6553]<=16'd57252;
ROM1[6554]<=16'd4743; ROM2[6554]<=16'd0; ROM3[6554]<=16'd23791; ROM4[6554]<=16'd57267;
ROM1[6555]<=16'd4763; ROM2[6555]<=16'd0; ROM3[6555]<=16'd23788; ROM4[6555]<=16'd57278;
ROM1[6556]<=16'd4786; ROM2[6556]<=16'd0; ROM3[6556]<=16'd23774; ROM4[6556]<=16'd57273;
ROM1[6557]<=16'd4815; ROM2[6557]<=16'd0; ROM3[6557]<=16'd23766; ROM4[6557]<=16'd57276;
ROM1[6558]<=16'd4816; ROM2[6558]<=16'd0; ROM3[6558]<=16'd23770; ROM4[6558]<=16'd57280;
ROM1[6559]<=16'd4808; ROM2[6559]<=16'd0; ROM3[6559]<=16'd23788; ROM4[6559]<=16'd57291;
ROM1[6560]<=16'd4799; ROM2[6560]<=16'd0; ROM3[6560]<=16'd23799; ROM4[6560]<=16'd57300;
ROM1[6561]<=16'd4777; ROM2[6561]<=16'd0; ROM3[6561]<=16'd23797; ROM4[6561]<=16'd57294;
ROM1[6562]<=16'd4765; ROM2[6562]<=16'd0; ROM3[6562]<=16'd23800; ROM4[6562]<=16'd57292;
ROM1[6563]<=16'd4770; ROM2[6563]<=16'd0; ROM3[6563]<=16'd23798; ROM4[6563]<=16'd57286;
ROM1[6564]<=16'd4787; ROM2[6564]<=16'd0; ROM3[6564]<=16'd23784; ROM4[6564]<=16'd57276;
ROM1[6565]<=16'd4815; ROM2[6565]<=16'd0; ROM3[6565]<=16'd23773; ROM4[6565]<=16'd57277;
ROM1[6566]<=16'd4822; ROM2[6566]<=16'd0; ROM3[6566]<=16'd23775; ROM4[6566]<=16'd57281;
ROM1[6567]<=16'd4822; ROM2[6567]<=16'd0; ROM3[6567]<=16'd23792; ROM4[6567]<=16'd57293;
ROM1[6568]<=16'd4814; ROM2[6568]<=16'd0; ROM3[6568]<=16'd23806; ROM4[6568]<=16'd57303;
ROM1[6569]<=16'd4788; ROM2[6569]<=16'd0; ROM3[6569]<=16'd23803; ROM4[6569]<=16'd57289;
ROM1[6570]<=16'd4759; ROM2[6570]<=16'd0; ROM3[6570]<=16'd23800; ROM4[6570]<=16'd57277;
ROM1[6571]<=16'd4761; ROM2[6571]<=16'd0; ROM3[6571]<=16'd23809; ROM4[6571]<=16'd57285;
ROM1[6572]<=16'd4791; ROM2[6572]<=16'd0; ROM3[6572]<=16'd23812; ROM4[6572]<=16'd57293;
ROM1[6573]<=16'd4808; ROM2[6573]<=16'd0; ROM3[6573]<=16'd23786; ROM4[6573]<=16'd57279;
ROM1[6574]<=16'd4816; ROM2[6574]<=16'd0; ROM3[6574]<=16'd23774; ROM4[6574]<=16'd57275;
ROM1[6575]<=16'd4792; ROM2[6575]<=16'd0; ROM3[6575]<=16'd23765; ROM4[6575]<=16'd57260;
ROM1[6576]<=16'd4767; ROM2[6576]<=16'd0; ROM3[6576]<=16'd23768; ROM4[6576]<=16'd57255;
ROM1[6577]<=16'd4767; ROM2[6577]<=16'd0; ROM3[6577]<=16'd23790; ROM4[6577]<=16'd57274;
ROM1[6578]<=16'd4757; ROM2[6578]<=16'd0; ROM3[6578]<=16'd23796; ROM4[6578]<=16'd57276;
ROM1[6579]<=16'd4742; ROM2[6579]<=16'd0; ROM3[6579]<=16'd23789; ROM4[6579]<=16'd57267;
ROM1[6580]<=16'd4741; ROM2[6580]<=16'd0; ROM3[6580]<=16'd23775; ROM4[6580]<=16'd57257;
ROM1[6581]<=16'd4775; ROM2[6581]<=16'd0; ROM3[6581]<=16'd23761; ROM4[6581]<=16'd57254;
ROM1[6582]<=16'd4809; ROM2[6582]<=16'd0; ROM3[6582]<=16'd23758; ROM4[6582]<=16'd57256;
ROM1[6583]<=16'd4806; ROM2[6583]<=16'd0; ROM3[6583]<=16'd23765; ROM4[6583]<=16'd57259;
ROM1[6584]<=16'd4791; ROM2[6584]<=16'd0; ROM3[6584]<=16'd23777; ROM4[6584]<=16'd57263;
ROM1[6585]<=16'd4790; ROM2[6585]<=16'd0; ROM3[6585]<=16'd23800; ROM4[6585]<=16'd57280;
ROM1[6586]<=16'd4770; ROM2[6586]<=16'd0; ROM3[6586]<=16'd23798; ROM4[6586]<=16'd57278;
ROM1[6587]<=16'd4745; ROM2[6587]<=16'd0; ROM3[6587]<=16'd23783; ROM4[6587]<=16'd57263;
ROM1[6588]<=16'd4752; ROM2[6588]<=16'd0; ROM3[6588]<=16'd23781; ROM4[6588]<=16'd57263;
ROM1[6589]<=16'd4767; ROM2[6589]<=16'd0; ROM3[6589]<=16'd23763; ROM4[6589]<=16'd57254;
ROM1[6590]<=16'd4800; ROM2[6590]<=16'd0; ROM3[6590]<=16'd23756; ROM4[6590]<=16'd57258;
ROM1[6591]<=16'd4807; ROM2[6591]<=16'd0; ROM3[6591]<=16'd23759; ROM4[6591]<=16'd57265;
ROM1[6592]<=16'd4779; ROM2[6592]<=16'd0; ROM3[6592]<=16'd23752; ROM4[6592]<=16'd57254;
ROM1[6593]<=16'd4754; ROM2[6593]<=16'd0; ROM3[6593]<=16'd23753; ROM4[6593]<=16'd57244;
ROM1[6594]<=16'd4735; ROM2[6594]<=16'd0; ROM3[6594]<=16'd23753; ROM4[6594]<=16'd57239;
ROM1[6595]<=16'd4725; ROM2[6595]<=16'd0; ROM3[6595]<=16'd23759; ROM4[6595]<=16'd57240;
ROM1[6596]<=16'd4745; ROM2[6596]<=16'd0; ROM3[6596]<=16'd23781; ROM4[6596]<=16'd57261;
ROM1[6597]<=16'd4785; ROM2[6597]<=16'd0; ROM3[6597]<=16'd23800; ROM4[6597]<=16'd57284;
ROM1[6598]<=16'd4815; ROM2[6598]<=16'd0; ROM3[6598]<=16'd23787; ROM4[6598]<=16'd57279;
ROM1[6599]<=16'd4809; ROM2[6599]<=16'd0; ROM3[6599]<=16'd23764; ROM4[6599]<=16'd57261;
ROM1[6600]<=16'd4781; ROM2[6600]<=16'd0; ROM3[6600]<=16'd23758; ROM4[6600]<=16'd57246;
ROM1[6601]<=16'd4757; ROM2[6601]<=16'd0; ROM3[6601]<=16'd23759; ROM4[6601]<=16'd57240;
ROM1[6602]<=16'd4764; ROM2[6602]<=16'd0; ROM3[6602]<=16'd23784; ROM4[6602]<=16'd57260;
ROM1[6603]<=16'd4782; ROM2[6603]<=16'd0; ROM3[6603]<=16'd23817; ROM4[6603]<=16'd57291;
ROM1[6604]<=16'd4780; ROM2[6604]<=16'd0; ROM3[6604]<=16'd23812; ROM4[6604]<=16'd57286;
ROM1[6605]<=16'd4772; ROM2[6605]<=16'd0; ROM3[6605]<=16'd23786; ROM4[6605]<=16'd57262;
ROM1[6606]<=16'd4794; ROM2[6606]<=16'd0; ROM3[6606]<=16'd23771; ROM4[6606]<=16'd57261;
ROM1[6607]<=16'd4814; ROM2[6607]<=16'd0; ROM3[6607]<=16'd23759; ROM4[6607]<=16'd57255;
ROM1[6608]<=16'd4807; ROM2[6608]<=16'd0; ROM3[6608]<=16'd23767; ROM4[6608]<=16'd57257;
ROM1[6609]<=16'd4796; ROM2[6609]<=16'd0; ROM3[6609]<=16'd23784; ROM4[6609]<=16'd57271;
ROM1[6610]<=16'd4781; ROM2[6610]<=16'd0; ROM3[6610]<=16'd23799; ROM4[6610]<=16'd57273;
ROM1[6611]<=16'd4766; ROM2[6611]<=16'd0; ROM3[6611]<=16'd23805; ROM4[6611]<=16'd57272;
ROM1[6612]<=16'd4754; ROM2[6612]<=16'd0; ROM3[6612]<=16'd23808; ROM4[6612]<=16'd57273;
ROM1[6613]<=16'd4763; ROM2[6613]<=16'd0; ROM3[6613]<=16'd23810; ROM4[6613]<=16'd57275;
ROM1[6614]<=16'd4793; ROM2[6614]<=16'd0; ROM3[6614]<=16'd23806; ROM4[6614]<=16'd57280;
ROM1[6615]<=16'd4824; ROM2[6615]<=16'd0; ROM3[6615]<=16'd23797; ROM4[6615]<=16'd57284;
ROM1[6616]<=16'd4823; ROM2[6616]<=16'd0; ROM3[6616]<=16'd23793; ROM4[6616]<=16'd57280;
ROM1[6617]<=16'd4809; ROM2[6617]<=16'd0; ROM3[6617]<=16'd23804; ROM4[6617]<=16'd57283;
ROM1[6618]<=16'd4788; ROM2[6618]<=16'd0; ROM3[6618]<=16'd23809; ROM4[6618]<=16'd57284;
ROM1[6619]<=16'd4793; ROM2[6619]<=16'd0; ROM3[6619]<=16'd23825; ROM4[6619]<=16'd57296;
ROM1[6620]<=16'd4790; ROM2[6620]<=16'd0; ROM3[6620]<=16'd23830; ROM4[6620]<=16'd57298;
ROM1[6621]<=16'd4774; ROM2[6621]<=16'd0; ROM3[6621]<=16'd23810; ROM4[6621]<=16'd57276;
ROM1[6622]<=16'd4777; ROM2[6622]<=16'd0; ROM3[6622]<=16'd23787; ROM4[6622]<=16'd57260;
ROM1[6623]<=16'd4809; ROM2[6623]<=16'd0; ROM3[6623]<=16'd23774; ROM4[6623]<=16'd57259;
ROM1[6624]<=16'd4838; ROM2[6624]<=16'd0; ROM3[6624]<=16'd23786; ROM4[6624]<=16'd57277;
ROM1[6625]<=16'd4845; ROM2[6625]<=16'd0; ROM3[6625]<=16'd23809; ROM4[6625]<=16'd57301;
ROM1[6626]<=16'd4828; ROM2[6626]<=16'd0; ROM3[6626]<=16'd23812; ROM4[6626]<=16'd57294;
ROM1[6627]<=16'd4797; ROM2[6627]<=16'd0; ROM3[6627]<=16'd23803; ROM4[6627]<=16'd57279;
ROM1[6628]<=16'd4779; ROM2[6628]<=16'd0; ROM3[6628]<=16'd23808; ROM4[6628]<=16'd57281;
ROM1[6629]<=16'd4761; ROM2[6629]<=16'd0; ROM3[6629]<=16'd23800; ROM4[6629]<=16'd57268;
ROM1[6630]<=16'd4771; ROM2[6630]<=16'd0; ROM3[6630]<=16'd23793; ROM4[6630]<=16'd57268;
ROM1[6631]<=16'd4805; ROM2[6631]<=16'd0; ROM3[6631]<=16'd23789; ROM4[6631]<=16'd57273;
ROM1[6632]<=16'd4825; ROM2[6632]<=16'd0; ROM3[6632]<=16'd23776; ROM4[6632]<=16'd57268;
ROM1[6633]<=16'd4822; ROM2[6633]<=16'd0; ROM3[6633]<=16'd23779; ROM4[6633]<=16'd57270;
ROM1[6634]<=16'd4800; ROM2[6634]<=16'd0; ROM3[6634]<=16'd23790; ROM4[6634]<=16'd57275;
ROM1[6635]<=16'd4782; ROM2[6635]<=16'd0; ROM3[6635]<=16'd23801; ROM4[6635]<=16'd57276;
ROM1[6636]<=16'd4772; ROM2[6636]<=16'd0; ROM3[6636]<=16'd23807; ROM4[6636]<=16'd57277;
ROM1[6637]<=16'd4755; ROM2[6637]<=16'd0; ROM3[6637]<=16'd23802; ROM4[6637]<=16'd57268;
ROM1[6638]<=16'd4769; ROM2[6638]<=16'd0; ROM3[6638]<=16'd23804; ROM4[6638]<=16'd57270;
ROM1[6639]<=16'd4800; ROM2[6639]<=16'd0; ROM3[6639]<=16'd23803; ROM4[6639]<=16'd57280;
ROM1[6640]<=16'd4819; ROM2[6640]<=16'd0; ROM3[6640]<=16'd23775; ROM4[6640]<=16'd57268;
ROM1[6641]<=16'd4827; ROM2[6641]<=16'd0; ROM3[6641]<=16'd23770; ROM4[6641]<=16'd57267;
ROM1[6642]<=16'd4811; ROM2[6642]<=16'd0; ROM3[6642]<=16'd23770; ROM4[6642]<=16'd57260;
ROM1[6643]<=16'd4773; ROM2[6643]<=16'd0; ROM3[6643]<=16'd23758; ROM4[6643]<=16'd57241;
ROM1[6644]<=16'd4762; ROM2[6644]<=16'd0; ROM3[6644]<=16'd23767; ROM4[6644]<=16'd57243;
ROM1[6645]<=16'd4759; ROM2[6645]<=16'd0; ROM3[6645]<=16'd23782; ROM4[6645]<=16'd57252;
ROM1[6646]<=16'd4766; ROM2[6646]<=16'd0; ROM3[6646]<=16'd23792; ROM4[6646]<=16'd57262;
ROM1[6647]<=16'd4804; ROM2[6647]<=16'd0; ROM3[6647]<=16'd23802; ROM4[6647]<=16'd57278;
ROM1[6648]<=16'd4833; ROM2[6648]<=16'd0; ROM3[6648]<=16'd23787; ROM4[6648]<=16'd57276;
ROM1[6649]<=16'd4846; ROM2[6649]<=16'd0; ROM3[6649]<=16'd23781; ROM4[6649]<=16'd57279;
ROM1[6650]<=16'd4831; ROM2[6650]<=16'd0; ROM3[6650]<=16'd23782; ROM4[6650]<=16'd57277;
ROM1[6651]<=16'd4796; ROM2[6651]<=16'd0; ROM3[6651]<=16'd23778; ROM4[6651]<=16'd57265;
ROM1[6652]<=16'd4785; ROM2[6652]<=16'd0; ROM3[6652]<=16'd23793; ROM4[6652]<=16'd57273;
ROM1[6653]<=16'd4771; ROM2[6653]<=16'd0; ROM3[6653]<=16'd23802; ROM4[6653]<=16'd57273;
ROM1[6654]<=16'd4766; ROM2[6654]<=16'd0; ROM3[6654]<=16'd23805; ROM4[6654]<=16'd57275;
ROM1[6655]<=16'd4783; ROM2[6655]<=16'd0; ROM3[6655]<=16'd23807; ROM4[6655]<=16'd57282;
ROM1[6656]<=16'd4810; ROM2[6656]<=16'd0; ROM3[6656]<=16'd23795; ROM4[6656]<=16'd57278;
ROM1[6657]<=16'd4829; ROM2[6657]<=16'd0; ROM3[6657]<=16'd23777; ROM4[6657]<=16'd57271;
ROM1[6658]<=16'd4818; ROM2[6658]<=16'd0; ROM3[6658]<=16'd23775; ROM4[6658]<=16'd57267;
ROM1[6659]<=16'd4801; ROM2[6659]<=16'd0; ROM3[6659]<=16'd23781; ROM4[6659]<=16'd57266;
ROM1[6660]<=16'd4785; ROM2[6660]<=16'd0; ROM3[6660]<=16'd23789; ROM4[6660]<=16'd57269;
ROM1[6661]<=16'd4776; ROM2[6661]<=16'd0; ROM3[6661]<=16'd23799; ROM4[6661]<=16'd57272;
ROM1[6662]<=16'd4771; ROM2[6662]<=16'd0; ROM3[6662]<=16'd23807; ROM4[6662]<=16'd57277;
ROM1[6663]<=16'd4784; ROM2[6663]<=16'd0; ROM3[6663]<=16'd23812; ROM4[6663]<=16'd57284;
ROM1[6664]<=16'd4806; ROM2[6664]<=16'd0; ROM3[6664]<=16'd23800; ROM4[6664]<=16'd57279;
ROM1[6665]<=16'd4822; ROM2[6665]<=16'd0; ROM3[6665]<=16'd23777; ROM4[6665]<=16'd57267;
ROM1[6666]<=16'd4824; ROM2[6666]<=16'd0; ROM3[6666]<=16'd23774; ROM4[6666]<=16'd57263;
ROM1[6667]<=16'd4815; ROM2[6667]<=16'd0; ROM3[6667]<=16'd23785; ROM4[6667]<=16'd57267;
ROM1[6668]<=16'd4803; ROM2[6668]<=16'd0; ROM3[6668]<=16'd23800; ROM4[6668]<=16'd57275;
ROM1[6669]<=16'd4797; ROM2[6669]<=16'd0; ROM3[6669]<=16'd23817; ROM4[6669]<=16'd57291;
ROM1[6670]<=16'd4769; ROM2[6670]<=16'd0; ROM3[6670]<=16'd23808; ROM4[6670]<=16'd57278;
ROM1[6671]<=16'd4752; ROM2[6671]<=16'd0; ROM3[6671]<=16'd23790; ROM4[6671]<=16'd57253;
ROM1[6672]<=16'd4769; ROM2[6672]<=16'd0; ROM3[6672]<=16'd23779; ROM4[6672]<=16'd57246;
ROM1[6673]<=16'd4800; ROM2[6673]<=16'd0; ROM3[6673]<=16'd23770; ROM4[6673]<=16'd57249;
ROM1[6674]<=16'd4814; ROM2[6674]<=16'd0; ROM3[6674]<=16'd23770; ROM4[6674]<=16'd57253;
ROM1[6675]<=16'd4798; ROM2[6675]<=16'd0; ROM3[6675]<=16'd23769; ROM4[6675]<=16'd57255;
ROM1[6676]<=16'd4786; ROM2[6676]<=16'd0; ROM3[6676]<=16'd23783; ROM4[6676]<=16'd57262;
ROM1[6677]<=16'd4782; ROM2[6677]<=16'd0; ROM3[6677]<=16'd23797; ROM4[6677]<=16'd57265;
ROM1[6678]<=16'd4763; ROM2[6678]<=16'd0; ROM3[6678]<=16'd23799; ROM4[6678]<=16'd57262;
ROM1[6679]<=16'd4754; ROM2[6679]<=16'd0; ROM3[6679]<=16'd23799; ROM4[6679]<=16'd57257;
ROM1[6680]<=16'd4778; ROM2[6680]<=16'd0; ROM3[6680]<=16'd23802; ROM4[6680]<=16'd57265;
ROM1[6681]<=16'd4801; ROM2[6681]<=16'd0; ROM3[6681]<=16'd23786; ROM4[6681]<=16'd57261;
ROM1[6682]<=16'd4810; ROM2[6682]<=16'd0; ROM3[6682]<=16'd23763; ROM4[6682]<=16'd57250;
ROM1[6683]<=16'd4802; ROM2[6683]<=16'd0; ROM3[6683]<=16'd23762; ROM4[6683]<=16'd57247;
ROM1[6684]<=16'd4782; ROM2[6684]<=16'd0; ROM3[6684]<=16'd23764; ROM4[6684]<=16'd57242;
ROM1[6685]<=16'd4769; ROM2[6685]<=16'd0; ROM3[6685]<=16'd23770; ROM4[6685]<=16'd57243;
ROM1[6686]<=16'd4763; ROM2[6686]<=16'd0; ROM3[6686]<=16'd23781; ROM4[6686]<=16'd57252;
ROM1[6687]<=16'd4749; ROM2[6687]<=16'd0; ROM3[6687]<=16'd23784; ROM4[6687]<=16'd57253;
ROM1[6688]<=16'd4743; ROM2[6688]<=16'd0; ROM3[6688]<=16'd23780; ROM4[6688]<=16'd57249;
ROM1[6689]<=16'd4762; ROM2[6689]<=16'd0; ROM3[6689]<=16'd23767; ROM4[6689]<=16'd57246;
ROM1[6690]<=16'd4799; ROM2[6690]<=16'd0; ROM3[6690]<=16'd23758; ROM4[6690]<=16'd57247;
ROM1[6691]<=16'd4806; ROM2[6691]<=16'd0; ROM3[6691]<=16'd23759; ROM4[6691]<=16'd57251;
ROM1[6692]<=16'd4787; ROM2[6692]<=16'd0; ROM3[6692]<=16'd23767; ROM4[6692]<=16'd57255;
ROM1[6693]<=16'd4771; ROM2[6693]<=16'd0; ROM3[6693]<=16'd23776; ROM4[6693]<=16'd57255;
ROM1[6694]<=16'd4764; ROM2[6694]<=16'd0; ROM3[6694]<=16'd23782; ROM4[6694]<=16'd57256;
ROM1[6695]<=16'd4746; ROM2[6695]<=16'd0; ROM3[6695]<=16'd23781; ROM4[6695]<=16'd57250;
ROM1[6696]<=16'd4738; ROM2[6696]<=16'd0; ROM3[6696]<=16'd23770; ROM4[6696]<=16'd57239;
ROM1[6697]<=16'd4752; ROM2[6697]<=16'd0; ROM3[6697]<=16'd23754; ROM4[6697]<=16'd57231;
ROM1[6698]<=16'd4778; ROM2[6698]<=16'd0; ROM3[6698]<=16'd23745; ROM4[6698]<=16'd57231;
ROM1[6699]<=16'd4802; ROM2[6699]<=16'd0; ROM3[6699]<=16'd23749; ROM4[6699]<=16'd57240;
ROM1[6700]<=16'd4802; ROM2[6700]<=16'd0; ROM3[6700]<=16'd23762; ROM4[6700]<=16'd57250;
ROM1[6701]<=16'd4784; ROM2[6701]<=16'd0; ROM3[6701]<=16'd23769; ROM4[6701]<=16'd57250;
ROM1[6702]<=16'd4776; ROM2[6702]<=16'd0; ROM3[6702]<=16'd23778; ROM4[6702]<=16'd57250;
ROM1[6703]<=16'd4759; ROM2[6703]<=16'd0; ROM3[6703]<=16'd23781; ROM4[6703]<=16'd57247;
ROM1[6704]<=16'd4730; ROM2[6704]<=16'd0; ROM3[6704]<=16'd23764; ROM4[6704]<=16'd57227;
ROM1[6705]<=16'd4740; ROM2[6705]<=16'd0; ROM3[6705]<=16'd23759; ROM4[6705]<=16'd57226;
ROM1[6706]<=16'd4773; ROM2[6706]<=16'd0; ROM3[6706]<=16'd23752; ROM4[6706]<=16'd57230;
ROM1[6707]<=16'd4801; ROM2[6707]<=16'd0; ROM3[6707]<=16'd23748; ROM4[6707]<=16'd57238;
ROM1[6708]<=16'd4803; ROM2[6708]<=16'd0; ROM3[6708]<=16'd23756; ROM4[6708]<=16'd57244;
ROM1[6709]<=16'd4780; ROM2[6709]<=16'd0; ROM3[6709]<=16'd23761; ROM4[6709]<=16'd57244;
ROM1[6710]<=16'd4770; ROM2[6710]<=16'd0; ROM3[6710]<=16'd23776; ROM4[6710]<=16'd57252;
ROM1[6711]<=16'd4770; ROM2[6711]<=16'd0; ROM3[6711]<=16'd23787; ROM4[6711]<=16'd57260;
ROM1[6712]<=16'd4763; ROM2[6712]<=16'd0; ROM3[6712]<=16'd23792; ROM4[6712]<=16'd57262;
ROM1[6713]<=16'd4775; ROM2[6713]<=16'd0; ROM3[6713]<=16'd23799; ROM4[6713]<=16'd57271;
ROM1[6714]<=16'd4799; ROM2[6714]<=16'd0; ROM3[6714]<=16'd23793; ROM4[6714]<=16'd57273;
ROM1[6715]<=16'd4821; ROM2[6715]<=16'd0; ROM3[6715]<=16'd23778; ROM4[6715]<=16'd57269;
ROM1[6716]<=16'd4827; ROM2[6716]<=16'd0; ROM3[6716]<=16'd23777; ROM4[6716]<=16'd57272;
ROM1[6717]<=16'd4818; ROM2[6717]<=16'd0; ROM3[6717]<=16'd23787; ROM4[6717]<=16'd57276;
ROM1[6718]<=16'd4806; ROM2[6718]<=16'd0; ROM3[6718]<=16'd23801; ROM4[6718]<=16'd57282;
ROM1[6719]<=16'd4797; ROM2[6719]<=16'd0; ROM3[6719]<=16'd23808; ROM4[6719]<=16'd57284;
ROM1[6720]<=16'd4775; ROM2[6720]<=16'd0; ROM3[6720]<=16'd23807; ROM4[6720]<=16'd57280;
ROM1[6721]<=16'd4770; ROM2[6721]<=16'd0; ROM3[6721]<=16'd23807; ROM4[6721]<=16'd57275;
ROM1[6722]<=16'd4796; ROM2[6722]<=16'd0; ROM3[6722]<=16'd23801; ROM4[6722]<=16'd57278;
ROM1[6723]<=16'd4828; ROM2[6723]<=16'd0; ROM3[6723]<=16'd23788; ROM4[6723]<=16'd57281;
ROM1[6724]<=16'd4850; ROM2[6724]<=16'd0; ROM3[6724]<=16'd23791; ROM4[6724]<=16'd57285;
ROM1[6725]<=16'd4861; ROM2[6725]<=16'd0; ROM3[6725]<=16'd23816; ROM4[6725]<=16'd57304;
ROM1[6726]<=16'd4841; ROM2[6726]<=16'd0; ROM3[6726]<=16'd23823; ROM4[6726]<=16'd57306;
ROM1[6727]<=16'd4799; ROM2[6727]<=16'd0; ROM3[6727]<=16'd23803; ROM4[6727]<=16'd57279;
ROM1[6728]<=16'd4771; ROM2[6728]<=16'd0; ROM3[6728]<=16'd23793; ROM4[6728]<=16'd57268;
ROM1[6729]<=16'd4761; ROM2[6729]<=16'd0; ROM3[6729]<=16'd23791; ROM4[6729]<=16'd57263;
ROM1[6730]<=16'd4766; ROM2[6730]<=16'd0; ROM3[6730]<=16'd23781; ROM4[6730]<=16'd57259;
ROM1[6731]<=16'd4800; ROM2[6731]<=16'd0; ROM3[6731]<=16'd23778; ROM4[6731]<=16'd57266;
ROM1[6732]<=16'd4824; ROM2[6732]<=16'd0; ROM3[6732]<=16'd23773; ROM4[6732]<=16'd57271;
ROM1[6733]<=16'd4803; ROM2[6733]<=16'd0; ROM3[6733]<=16'd23763; ROM4[6733]<=16'd57261;
ROM1[6734]<=16'd4784; ROM2[6734]<=16'd0; ROM3[6734]<=16'd23767; ROM4[6734]<=16'd57255;
ROM1[6735]<=16'd4781; ROM2[6735]<=16'd0; ROM3[6735]<=16'd23783; ROM4[6735]<=16'd57263;
ROM1[6736]<=16'd4786; ROM2[6736]<=16'd0; ROM3[6736]<=16'd23809; ROM4[6736]<=16'd57286;
ROM1[6737]<=16'd4780; ROM2[6737]<=16'd0; ROM3[6737]<=16'd23816; ROM4[6737]<=16'd57294;
ROM1[6738]<=16'd4776; ROM2[6738]<=16'd0; ROM3[6738]<=16'd23803; ROM4[6738]<=16'd57283;
ROM1[6739]<=16'd4795; ROM2[6739]<=16'd0; ROM3[6739]<=16'd23794; ROM4[6739]<=16'd57282;
ROM1[6740]<=16'd4823; ROM2[6740]<=16'd0; ROM3[6740]<=16'd23777; ROM4[6740]<=16'd57275;
ROM1[6741]<=16'd4827; ROM2[6741]<=16'd0; ROM3[6741]<=16'd23772; ROM4[6741]<=16'd57271;
ROM1[6742]<=16'd4813; ROM2[6742]<=16'd0; ROM3[6742]<=16'd23779; ROM4[6742]<=16'd57275;
ROM1[6743]<=16'd4801; ROM2[6743]<=16'd0; ROM3[6743]<=16'd23788; ROM4[6743]<=16'd57276;
ROM1[6744]<=16'd4799; ROM2[6744]<=16'd0; ROM3[6744]<=16'd23802; ROM4[6744]<=16'd57285;
ROM1[6745]<=16'd4809; ROM2[6745]<=16'd0; ROM3[6745]<=16'd23832; ROM4[6745]<=16'd57308;
ROM1[6746]<=16'd4815; ROM2[6746]<=16'd0; ROM3[6746]<=16'd23839; ROM4[6746]<=16'd57317;
ROM1[6747]<=16'd4816; ROM2[6747]<=16'd0; ROM3[6747]<=16'd23819; ROM4[6747]<=16'd57305;
ROM1[6748]<=16'd4830; ROM2[6748]<=16'd0; ROM3[6748]<=16'd23795; ROM4[6748]<=16'd57286;
ROM1[6749]<=16'd4819; ROM2[6749]<=16'd0; ROM3[6749]<=16'd23766; ROM4[6749]<=16'd57263;
ROM1[6750]<=16'd4801; ROM2[6750]<=16'd0; ROM3[6750]<=16'd23760; ROM4[6750]<=16'd57257;
ROM1[6751]<=16'd4796; ROM2[6751]<=16'd0; ROM3[6751]<=16'd23775; ROM4[6751]<=16'd57272;
ROM1[6752]<=16'd4788; ROM2[6752]<=16'd0; ROM3[6752]<=16'd23781; ROM4[6752]<=16'd57276;
ROM1[6753]<=16'd4768; ROM2[6753]<=16'd0; ROM3[6753]<=16'd23787; ROM4[6753]<=16'd57269;
ROM1[6754]<=16'd4759; ROM2[6754]<=16'd0; ROM3[6754]<=16'd23791; ROM4[6754]<=16'd57267;
ROM1[6755]<=16'd4769; ROM2[6755]<=16'd0; ROM3[6755]<=16'd23781; ROM4[6755]<=16'd57263;
ROM1[6756]<=16'd4784; ROM2[6756]<=16'd0; ROM3[6756]<=16'd23756; ROM4[6756]<=16'd57248;
ROM1[6757]<=16'd4802; ROM2[6757]<=16'd0; ROM3[6757]<=16'd23739; ROM4[6757]<=16'd57244;
ROM1[6758]<=16'd4800; ROM2[6758]<=16'd0; ROM3[6758]<=16'd23746; ROM4[6758]<=16'd57249;
ROM1[6759]<=16'd4787; ROM2[6759]<=16'd0; ROM3[6759]<=16'd23762; ROM4[6759]<=16'd57252;
ROM1[6760]<=16'd4776; ROM2[6760]<=16'd0; ROM3[6760]<=16'd23775; ROM4[6760]<=16'd57258;
ROM1[6761]<=16'd4765; ROM2[6761]<=16'd0; ROM3[6761]<=16'd23782; ROM4[6761]<=16'd57261;
ROM1[6762]<=16'd4760; ROM2[6762]<=16'd0; ROM3[6762]<=16'd23788; ROM4[6762]<=16'd57267;
ROM1[6763]<=16'd4766; ROM2[6763]<=16'd0; ROM3[6763]<=16'd23787; ROM4[6763]<=16'd57268;
ROM1[6764]<=16'd4793; ROM2[6764]<=16'd0; ROM3[6764]<=16'd23783; ROM4[6764]<=16'd57273;
ROM1[6765]<=16'd4832; ROM2[6765]<=16'd0; ROM3[6765]<=16'd23782; ROM4[6765]<=16'd57283;
ROM1[6766]<=16'd4833; ROM2[6766]<=16'd0; ROM3[6766]<=16'd23778; ROM4[6766]<=16'd57276;
ROM1[6767]<=16'd4820; ROM2[6767]<=16'd0; ROM3[6767]<=16'd23785; ROM4[6767]<=16'd57281;
ROM1[6768]<=16'd4799; ROM2[6768]<=16'd0; ROM3[6768]<=16'd23789; ROM4[6768]<=16'd57278;
ROM1[6769]<=16'd4776; ROM2[6769]<=16'd0; ROM3[6769]<=16'd23785; ROM4[6769]<=16'd57271;
ROM1[6770]<=16'd4764; ROM2[6770]<=16'd0; ROM3[6770]<=16'd23792; ROM4[6770]<=16'd57277;
ROM1[6771]<=16'd4770; ROM2[6771]<=16'd0; ROM3[6771]<=16'd23804; ROM4[6771]<=16'd57282;
ROM1[6772]<=16'd4794; ROM2[6772]<=16'd0; ROM3[6772]<=16'd23804; ROM4[6772]<=16'd57284;
ROM1[6773]<=16'd4819; ROM2[6773]<=16'd0; ROM3[6773]<=16'd23784; ROM4[6773]<=16'd57278;
ROM1[6774]<=16'd4818; ROM2[6774]<=16'd0; ROM3[6774]<=16'd23770; ROM4[6774]<=16'd57268;
ROM1[6775]<=16'd4806; ROM2[6775]<=16'd0; ROM3[6775]<=16'd23776; ROM4[6775]<=16'd57271;
ROM1[6776]<=16'd4799; ROM2[6776]<=16'd0; ROM3[6776]<=16'd23791; ROM4[6776]<=16'd57286;
ROM1[6777]<=16'd4789; ROM2[6777]<=16'd0; ROM3[6777]<=16'd23800; ROM4[6777]<=16'd57287;
ROM1[6778]<=16'd4770; ROM2[6778]<=16'd0; ROM3[6778]<=16'd23805; ROM4[6778]<=16'd57284;
ROM1[6779]<=16'd4757; ROM2[6779]<=16'd0; ROM3[6779]<=16'd23806; ROM4[6779]<=16'd57285;
ROM1[6780]<=16'd4761; ROM2[6780]<=16'd0; ROM3[6780]<=16'd23796; ROM4[6780]<=16'd57279;
ROM1[6781]<=16'd4797; ROM2[6781]<=16'd0; ROM3[6781]<=16'd23785; ROM4[6781]<=16'd57283;
ROM1[6782]<=16'd4825; ROM2[6782]<=16'd0; ROM3[6782]<=16'd23778; ROM4[6782]<=16'd57289;
ROM1[6783]<=16'd4816; ROM2[6783]<=16'd0; ROM3[6783]<=16'd23777; ROM4[6783]<=16'd57288;
ROM1[6784]<=16'd4800; ROM2[6784]<=16'd0; ROM3[6784]<=16'd23784; ROM4[6784]<=16'd57290;
ROM1[6785]<=16'd4790; ROM2[6785]<=16'd0; ROM3[6785]<=16'd23799; ROM4[6785]<=16'd57298;
ROM1[6786]<=16'd4787; ROM2[6786]<=16'd0; ROM3[6786]<=16'd23808; ROM4[6786]<=16'd57301;
ROM1[6787]<=16'd4776; ROM2[6787]<=16'd0; ROM3[6787]<=16'd23809; ROM4[6787]<=16'd57296;
ROM1[6788]<=16'd4775; ROM2[6788]<=16'd0; ROM3[6788]<=16'd23800; ROM4[6788]<=16'd57294;
ROM1[6789]<=16'd4811; ROM2[6789]<=16'd0; ROM3[6789]<=16'd23806; ROM4[6789]<=16'd57308;
ROM1[6790]<=16'd4878; ROM2[6790]<=16'd0; ROM3[6790]<=16'd23836; ROM4[6790]<=16'd57346;
ROM1[6791]<=16'd4875; ROM2[6791]<=16'd0; ROM3[6791]<=16'd23829; ROM4[6791]<=16'd57338;
ROM1[6792]<=16'd4830; ROM2[6792]<=16'd0; ROM3[6792]<=16'd23803; ROM4[6792]<=16'd57305;
ROM1[6793]<=16'd4796; ROM2[6793]<=16'd0; ROM3[6793]<=16'd23794; ROM4[6793]<=16'd57287;
ROM1[6794]<=16'd4765; ROM2[6794]<=16'd0; ROM3[6794]<=16'd23785; ROM4[6794]<=16'd57270;
ROM1[6795]<=16'd4749; ROM2[6795]<=16'd0; ROM3[6795]<=16'd23790; ROM4[6795]<=16'd57263;
ROM1[6796]<=16'd4760; ROM2[6796]<=16'd0; ROM3[6796]<=16'd23801; ROM4[6796]<=16'd57273;
ROM1[6797]<=16'd4782; ROM2[6797]<=16'd0; ROM3[6797]<=16'd23796; ROM4[6797]<=16'd57274;
ROM1[6798]<=16'd4804; ROM2[6798]<=16'd0; ROM3[6798]<=16'd23778; ROM4[6798]<=16'd57267;
ROM1[6799]<=16'd4826; ROM2[6799]<=16'd0; ROM3[6799]<=16'd23781; ROM4[6799]<=16'd57278;
ROM1[6800]<=16'd4824; ROM2[6800]<=16'd0; ROM3[6800]<=16'd23792; ROM4[6800]<=16'd57286;
ROM1[6801]<=16'd4791; ROM2[6801]<=16'd0; ROM3[6801]<=16'd23788; ROM4[6801]<=16'd57273;
ROM1[6802]<=16'd4772; ROM2[6802]<=16'd0; ROM3[6802]<=16'd23784; ROM4[6802]<=16'd57268;
ROM1[6803]<=16'd4761; ROM2[6803]<=16'd0; ROM3[6803]<=16'd23789; ROM4[6803]<=16'd57269;
ROM1[6804]<=16'd4756; ROM2[6804]<=16'd0; ROM3[6804]<=16'd23794; ROM4[6804]<=16'd57270;
ROM1[6805]<=16'd4767; ROM2[6805]<=16'd0; ROM3[6805]<=16'd23787; ROM4[6805]<=16'd57266;
ROM1[6806]<=16'd4789; ROM2[6806]<=16'd0; ROM3[6806]<=16'd23765; ROM4[6806]<=16'd57254;
ROM1[6807]<=16'd4809; ROM2[6807]<=16'd0; ROM3[6807]<=16'd23752; ROM4[6807]<=16'd57253;
ROM1[6808]<=16'd4811; ROM2[6808]<=16'd0; ROM3[6808]<=16'd23760; ROM4[6808]<=16'd57259;
ROM1[6809]<=16'd4806; ROM2[6809]<=16'd0; ROM3[6809]<=16'd23776; ROM4[6809]<=16'd57269;
ROM1[6810]<=16'd4785; ROM2[6810]<=16'd0; ROM3[6810]<=16'd23780; ROM4[6810]<=16'd57269;
ROM1[6811]<=16'd4764; ROM2[6811]<=16'd0; ROM3[6811]<=16'd23777; ROM4[6811]<=16'd57262;
ROM1[6812]<=16'd4760; ROM2[6812]<=16'd0; ROM3[6812]<=16'd23786; ROM4[6812]<=16'd57268;
ROM1[6813]<=16'd4765; ROM2[6813]<=16'd0; ROM3[6813]<=16'd23783; ROM4[6813]<=16'd57270;
ROM1[6814]<=16'd4787; ROM2[6814]<=16'd0; ROM3[6814]<=16'd23767; ROM4[6814]<=16'd57260;
ROM1[6815]<=16'd4820; ROM2[6815]<=16'd0; ROM3[6815]<=16'd23758; ROM4[6815]<=16'd57261;
ROM1[6816]<=16'd4824; ROM2[6816]<=16'd0; ROM3[6816]<=16'd23764; ROM4[6816]<=16'd57266;
ROM1[6817]<=16'd4810; ROM2[6817]<=16'd0; ROM3[6817]<=16'd23774; ROM4[6817]<=16'd57269;
ROM1[6818]<=16'd4794; ROM2[6818]<=16'd0; ROM3[6818]<=16'd23784; ROM4[6818]<=16'd57273;
ROM1[6819]<=16'd4781; ROM2[6819]<=16'd0; ROM3[6819]<=16'd23789; ROM4[6819]<=16'd57271;
ROM1[6820]<=16'd4769; ROM2[6820]<=16'd0; ROM3[6820]<=16'd23791; ROM4[6820]<=16'd57273;
ROM1[6821]<=16'd4795; ROM2[6821]<=16'd0; ROM3[6821]<=16'd23819; ROM4[6821]<=16'd57297;
ROM1[6822]<=16'd4822; ROM2[6822]<=16'd0; ROM3[6822]<=16'd23825; ROM4[6822]<=16'd57305;
ROM1[6823]<=16'd4831; ROM2[6823]<=16'd0; ROM3[6823]<=16'd23789; ROM4[6823]<=16'd57289;
ROM1[6824]<=16'd4853; ROM2[6824]<=16'd0; ROM3[6824]<=16'd23791; ROM4[6824]<=16'd57298;
ROM1[6825]<=16'd4822; ROM2[6825]<=16'd0; ROM3[6825]<=16'd23774; ROM4[6825]<=16'd57278;
ROM1[6826]<=16'd4784; ROM2[6826]<=16'd0; ROM3[6826]<=16'd23760; ROM4[6826]<=16'd57259;
ROM1[6827]<=16'd4781; ROM2[6827]<=16'd0; ROM3[6827]<=16'd23775; ROM4[6827]<=16'd57269;
ROM1[6828]<=16'd4754; ROM2[6828]<=16'd0; ROM3[6828]<=16'd23771; ROM4[6828]<=16'd57260;
ROM1[6829]<=16'd4740; ROM2[6829]<=16'd0; ROM3[6829]<=16'd23770; ROM4[6829]<=16'd57252;
ROM1[6830]<=16'd4758; ROM2[6830]<=16'd0; ROM3[6830]<=16'd23766; ROM4[6830]<=16'd57256;
ROM1[6831]<=16'd4791; ROM2[6831]<=16'd0; ROM3[6831]<=16'd23759; ROM4[6831]<=16'd57256;
ROM1[6832]<=16'd4806; ROM2[6832]<=16'd0; ROM3[6832]<=16'd23747; ROM4[6832]<=16'd57247;
ROM1[6833]<=16'd4796; ROM2[6833]<=16'd0; ROM3[6833]<=16'd23744; ROM4[6833]<=16'd57244;
ROM1[6834]<=16'd4790; ROM2[6834]<=16'd0; ROM3[6834]<=16'd23759; ROM4[6834]<=16'd57251;
ROM1[6835]<=16'd4790; ROM2[6835]<=16'd0; ROM3[6835]<=16'd23777; ROM4[6835]<=16'd57266;
ROM1[6836]<=16'd4786; ROM2[6836]<=16'd0; ROM3[6836]<=16'd23788; ROM4[6836]<=16'd57278;
ROM1[6837]<=16'd4780; ROM2[6837]<=16'd0; ROM3[6837]<=16'd23798; ROM4[6837]<=16'd57282;
ROM1[6838]<=16'd4792; ROM2[6838]<=16'd0; ROM3[6838]<=16'd23803; ROM4[6838]<=16'd57290;
ROM1[6839]<=16'd4820; ROM2[6839]<=16'd0; ROM3[6839]<=16'd23802; ROM4[6839]<=16'd57295;
ROM1[6840]<=16'd4842; ROM2[6840]<=16'd0; ROM3[6840]<=16'd23782; ROM4[6840]<=16'd57285;
ROM1[6841]<=16'd4837; ROM2[6841]<=16'd0; ROM3[6841]<=16'd23768; ROM4[6841]<=16'd57276;
ROM1[6842]<=16'd4817; ROM2[6842]<=16'd0; ROM3[6842]<=16'd23775; ROM4[6842]<=16'd57278;
ROM1[6843]<=16'd4796; ROM2[6843]<=16'd0; ROM3[6843]<=16'd23781; ROM4[6843]<=16'd57274;
ROM1[6844]<=16'd4787; ROM2[6844]<=16'd0; ROM3[6844]<=16'd23788; ROM4[6844]<=16'd57279;
ROM1[6845]<=16'd4776; ROM2[6845]<=16'd0; ROM3[6845]<=16'd23791; ROM4[6845]<=16'd57283;
ROM1[6846]<=16'd4775; ROM2[6846]<=16'd0; ROM3[6846]<=16'd23790; ROM4[6846]<=16'd57284;
ROM1[6847]<=16'd4792; ROM2[6847]<=16'd0; ROM3[6847]<=16'd23784; ROM4[6847]<=16'd57284;
ROM1[6848]<=16'd4823; ROM2[6848]<=16'd0; ROM3[6848]<=16'd23771; ROM4[6848]<=16'd57282;
ROM1[6849]<=16'd4827; ROM2[6849]<=16'd0; ROM3[6849]<=16'd23763; ROM4[6849]<=16'd57275;
ROM1[6850]<=16'd4812; ROM2[6850]<=16'd0; ROM3[6850]<=16'd23767; ROM4[6850]<=16'd57275;
ROM1[6851]<=16'd4802; ROM2[6851]<=16'd0; ROM3[6851]<=16'd23778; ROM4[6851]<=16'd57278;
ROM1[6852]<=16'd4795; ROM2[6852]<=16'd0; ROM3[6852]<=16'd23792; ROM4[6852]<=16'd57286;
ROM1[6853]<=16'd4786; ROM2[6853]<=16'd0; ROM3[6853]<=16'd23802; ROM4[6853]<=16'd57291;
ROM1[6854]<=16'd4762; ROM2[6854]<=16'd0; ROM3[6854]<=16'd23782; ROM4[6854]<=16'd57270;
ROM1[6855]<=16'd4755; ROM2[6855]<=16'd0; ROM3[6855]<=16'd23764; ROM4[6855]<=16'd57255;
ROM1[6856]<=16'd4781; ROM2[6856]<=16'd0; ROM3[6856]<=16'd23747; ROM4[6856]<=16'd57249;
ROM1[6857]<=16'd4809; ROM2[6857]<=16'd0; ROM3[6857]<=16'd23741; ROM4[6857]<=16'd57252;
ROM1[6858]<=16'd4826; ROM2[6858]<=16'd0; ROM3[6858]<=16'd23765; ROM4[6858]<=16'd57273;
ROM1[6859]<=16'd4807; ROM2[6859]<=16'd0; ROM3[6859]<=16'd23771; ROM4[6859]<=16'd57271;
ROM1[6860]<=16'd4774; ROM2[6860]<=16'd0; ROM3[6860]<=16'd23765; ROM4[6860]<=16'd57259;
ROM1[6861]<=16'd4757; ROM2[6861]<=16'd0; ROM3[6861]<=16'd23770; ROM4[6861]<=16'd57263;
ROM1[6862]<=16'd4734; ROM2[6862]<=16'd0; ROM3[6862]<=16'd23757; ROM4[6862]<=16'd57249;
ROM1[6863]<=16'd4739; ROM2[6863]<=16'd0; ROM3[6863]<=16'd23748; ROM4[6863]<=16'd57242;
ROM1[6864]<=16'd4768; ROM2[6864]<=16'd0; ROM3[6864]<=16'd23745; ROM4[6864]<=16'd57247;
ROM1[6865]<=16'd4801; ROM2[6865]<=16'd0; ROM3[6865]<=16'd23739; ROM4[6865]<=16'd57248;
ROM1[6866]<=16'd4823; ROM2[6866]<=16'd0; ROM3[6866]<=16'd23757; ROM4[6866]<=16'd57270;
ROM1[6867]<=16'd4805; ROM2[6867]<=16'd0; ROM3[6867]<=16'd23760; ROM4[6867]<=16'd57268;
ROM1[6868]<=16'd4776; ROM2[6868]<=16'd0; ROM3[6868]<=16'd23752; ROM4[6868]<=16'd57250;
ROM1[6869]<=16'd4758; ROM2[6869]<=16'd0; ROM3[6869]<=16'd23752; ROM4[6869]<=16'd57246;
ROM1[6870]<=16'd4740; ROM2[6870]<=16'd0; ROM3[6870]<=16'd23759; ROM4[6870]<=16'd57247;
ROM1[6871]<=16'd4749; ROM2[6871]<=16'd0; ROM3[6871]<=16'd23768; ROM4[6871]<=16'd57256;
ROM1[6872]<=16'd4785; ROM2[6872]<=16'd0; ROM3[6872]<=16'd23775; ROM4[6872]<=16'd57271;
ROM1[6873]<=16'd4835; ROM2[6873]<=16'd0; ROM3[6873]<=16'd23780; ROM4[6873]<=16'd57286;
ROM1[6874]<=16'd4858; ROM2[6874]<=16'd0; ROM3[6874]<=16'd23783; ROM4[6874]<=16'd57292;
ROM1[6875]<=16'd4856; ROM2[6875]<=16'd0; ROM3[6875]<=16'd23797; ROM4[6875]<=16'd57305;
ROM1[6876]<=16'd4825; ROM2[6876]<=16'd0; ROM3[6876]<=16'd23790; ROM4[6876]<=16'd57294;
ROM1[6877]<=16'd4800; ROM2[6877]<=16'd0; ROM3[6877]<=16'd23781; ROM4[6877]<=16'd57276;
ROM1[6878]<=16'd4789; ROM2[6878]<=16'd0; ROM3[6878]<=16'd23786; ROM4[6878]<=16'd57276;
ROM1[6879]<=16'd4776; ROM2[6879]<=16'd0; ROM3[6879]<=16'd23782; ROM4[6879]<=16'd57268;
ROM1[6880]<=16'd4798; ROM2[6880]<=16'd0; ROM3[6880]<=16'd23790; ROM4[6880]<=16'd57274;
ROM1[6881]<=16'd4838; ROM2[6881]<=16'd0; ROM3[6881]<=16'd23788; ROM4[6881]<=16'd57285;
ROM1[6882]<=16'd4835; ROM2[6882]<=16'd0; ROM3[6882]<=16'd23753; ROM4[6882]<=16'd57261;
ROM1[6883]<=16'd4812; ROM2[6883]<=16'd0; ROM3[6883]<=16'd23732; ROM4[6883]<=16'd57243;
ROM1[6884]<=16'd4797; ROM2[6884]<=16'd0; ROM3[6884]<=16'd23739; ROM4[6884]<=16'd57249;
ROM1[6885]<=16'd4771; ROM2[6885]<=16'd0; ROM3[6885]<=16'd23736; ROM4[6885]<=16'd57241;
ROM1[6886]<=16'd4760; ROM2[6886]<=16'd0; ROM3[6886]<=16'd23744; ROM4[6886]<=16'd57244;
ROM1[6887]<=16'd4760; ROM2[6887]<=16'd0; ROM3[6887]<=16'd23759; ROM4[6887]<=16'd57252;
ROM1[6888]<=16'd4766; ROM2[6888]<=16'd0; ROM3[6888]<=16'd23755; ROM4[6888]<=16'd57250;
ROM1[6889]<=16'd4801; ROM2[6889]<=16'd0; ROM3[6889]<=16'd23751; ROM4[6889]<=16'd57256;
ROM1[6890]<=16'd4832; ROM2[6890]<=16'd0; ROM3[6890]<=16'd23740; ROM4[6890]<=16'd57258;
ROM1[6891]<=16'd4822; ROM2[6891]<=16'd0; ROM3[6891]<=16'd23730; ROM4[6891]<=16'd57251;
ROM1[6892]<=16'd4803; ROM2[6892]<=16'd0; ROM3[6892]<=16'd23737; ROM4[6892]<=16'd57249;
ROM1[6893]<=16'd4789; ROM2[6893]<=16'd0; ROM3[6893]<=16'd23754; ROM4[6893]<=16'd57259;
ROM1[6894]<=16'd4798; ROM2[6894]<=16'd0; ROM3[6894]<=16'd23784; ROM4[6894]<=16'd57283;
ROM1[6895]<=16'd4819; ROM2[6895]<=16'd0; ROM3[6895]<=16'd23817; ROM4[6895]<=16'd57312;
ROM1[6896]<=16'd4813; ROM2[6896]<=16'd0; ROM3[6896]<=16'd23806; ROM4[6896]<=16'd57306;
ROM1[6897]<=16'd4802; ROM2[6897]<=16'd0; ROM3[6897]<=16'd23769; ROM4[6897]<=16'd57277;
ROM1[6898]<=16'd4823; ROM2[6898]<=16'd0; ROM3[6898]<=16'd23751; ROM4[6898]<=16'd57269;
ROM1[6899]<=16'd4830; ROM2[6899]<=16'd0; ROM3[6899]<=16'd23739; ROM4[6899]<=16'd57266;
ROM1[6900]<=16'd4824; ROM2[6900]<=16'd0; ROM3[6900]<=16'd23753; ROM4[6900]<=16'd57272;
ROM1[6901]<=16'd4820; ROM2[6901]<=16'd0; ROM3[6901]<=16'd23776; ROM4[6901]<=16'd57288;
ROM1[6902]<=16'd4810; ROM2[6902]<=16'd0; ROM3[6902]<=16'd23782; ROM4[6902]<=16'd57293;
ROM1[6903]<=16'd4795; ROM2[6903]<=16'd0; ROM3[6903]<=16'd23794; ROM4[6903]<=16'd57295;
ROM1[6904]<=16'd4794; ROM2[6904]<=16'd0; ROM3[6904]<=16'd23799; ROM4[6904]<=16'd57300;
ROM1[6905]<=16'd4802; ROM2[6905]<=16'd0; ROM3[6905]<=16'd23789; ROM4[6905]<=16'd57294;
ROM1[6906]<=16'd4821; ROM2[6906]<=16'd0; ROM3[6906]<=16'd23773; ROM4[6906]<=16'd57284;
ROM1[6907]<=16'd4840; ROM2[6907]<=16'd0; ROM3[6907]<=16'd23763; ROM4[6907]<=16'd57282;
ROM1[6908]<=16'd4830; ROM2[6908]<=16'd0; ROM3[6908]<=16'd23760; ROM4[6908]<=16'd57280;
ROM1[6909]<=16'd4812; ROM2[6909]<=16'd0; ROM3[6909]<=16'd23765; ROM4[6909]<=16'd57281;
ROM1[6910]<=16'd4794; ROM2[6910]<=16'd0; ROM3[6910]<=16'd23768; ROM4[6910]<=16'd57275;
ROM1[6911]<=16'd4773; ROM2[6911]<=16'd0; ROM3[6911]<=16'd23766; ROM4[6911]<=16'd57266;
ROM1[6912]<=16'd4761; ROM2[6912]<=16'd0; ROM3[6912]<=16'd23770; ROM4[6912]<=16'd57265;
ROM1[6913]<=16'd4770; ROM2[6913]<=16'd0; ROM3[6913]<=16'd23768; ROM4[6913]<=16'd57263;
ROM1[6914]<=16'd4793; ROM2[6914]<=16'd0; ROM3[6914]<=16'd23747; ROM4[6914]<=16'd57255;
ROM1[6915]<=16'd4814; ROM2[6915]<=16'd0; ROM3[6915]<=16'd23726; ROM4[6915]<=16'd57244;
ROM1[6916]<=16'd4810; ROM2[6916]<=16'd0; ROM3[6916]<=16'd23717; ROM4[6916]<=16'd57240;
ROM1[6917]<=16'd4792; ROM2[6917]<=16'd0; ROM3[6917]<=16'd23720; ROM4[6917]<=16'd57239;
ROM1[6918]<=16'd4782; ROM2[6918]<=16'd0; ROM3[6918]<=16'd23736; ROM4[6918]<=16'd57250;
ROM1[6919]<=16'd4780; ROM2[6919]<=16'd0; ROM3[6919]<=16'd23754; ROM4[6919]<=16'd57267;
ROM1[6920]<=16'd4769; ROM2[6920]<=16'd0; ROM3[6920]<=16'd23764; ROM4[6920]<=16'd57270;
ROM1[6921]<=16'd4769; ROM2[6921]<=16'd0; ROM3[6921]<=16'd23768; ROM4[6921]<=16'd57272;
ROM1[6922]<=16'd4792; ROM2[6922]<=16'd0; ROM3[6922]<=16'd23767; ROM4[6922]<=16'd57279;
ROM1[6923]<=16'd4815; ROM2[6923]<=16'd0; ROM3[6923]<=16'd23745; ROM4[6923]<=16'd57272;
ROM1[6924]<=16'd4823; ROM2[6924]<=16'd0; ROM3[6924]<=16'd23732; ROM4[6924]<=16'd57264;
ROM1[6925]<=16'd4804; ROM2[6925]<=16'd0; ROM3[6925]<=16'd23735; ROM4[6925]<=16'd57259;
ROM1[6926]<=16'd4776; ROM2[6926]<=16'd0; ROM3[6926]<=16'd23739; ROM4[6926]<=16'd57253;
ROM1[6927]<=16'd4774; ROM2[6927]<=16'd0; ROM3[6927]<=16'd23761; ROM4[6927]<=16'd57267;
ROM1[6928]<=16'd4757; ROM2[6928]<=16'd0; ROM3[6928]<=16'd23775; ROM4[6928]<=16'd57275;
ROM1[6929]<=16'd4744; ROM2[6929]<=16'd0; ROM3[6929]<=16'd23769; ROM4[6929]<=16'd57265;
ROM1[6930]<=16'd4761; ROM2[6930]<=16'd0; ROM3[6930]<=16'd23767; ROM4[6930]<=16'd57267;
ROM1[6931]<=16'd4796; ROM2[6931]<=16'd0; ROM3[6931]<=16'd23761; ROM4[6931]<=16'd57273;
ROM1[6932]<=16'd4827; ROM2[6932]<=16'd0; ROM3[6932]<=16'd23759; ROM4[6932]<=16'd57279;
ROM1[6933]<=16'd4826; ROM2[6933]<=16'd0; ROM3[6933]<=16'd23765; ROM4[6933]<=16'd57289;
ROM1[6934]<=16'd4808; ROM2[6934]<=16'd0; ROM3[6934]<=16'd23772; ROM4[6934]<=16'd57285;
ROM1[6935]<=16'd4784; ROM2[6935]<=16'd0; ROM3[6935]<=16'd23767; ROM4[6935]<=16'd57272;
ROM1[6936]<=16'd4766; ROM2[6936]<=16'd0; ROM3[6936]<=16'd23766; ROM4[6936]<=16'd57269;
ROM1[6937]<=16'd4752; ROM2[6937]<=16'd0; ROM3[6937]<=16'd23765; ROM4[6937]<=16'd57264;
ROM1[6938]<=16'd4756; ROM2[6938]<=16'd0; ROM3[6938]<=16'd23757; ROM4[6938]<=16'd57263;
ROM1[6939]<=16'd4781; ROM2[6939]<=16'd0; ROM3[6939]<=16'd23746; ROM4[6939]<=16'd57265;
ROM1[6940]<=16'd4809; ROM2[6940]<=16'd0; ROM3[6940]<=16'd23733; ROM4[6940]<=16'd57266;
ROM1[6941]<=16'd4822; ROM2[6941]<=16'd0; ROM3[6941]<=16'd23738; ROM4[6941]<=16'd57274;
ROM1[6942]<=16'd4812; ROM2[6942]<=16'd0; ROM3[6942]<=16'd23749; ROM4[6942]<=16'd57280;
ROM1[6943]<=16'd4787; ROM2[6943]<=16'd0; ROM3[6943]<=16'd23753; ROM4[6943]<=16'd57274;
ROM1[6944]<=16'd4766; ROM2[6944]<=16'd0; ROM3[6944]<=16'd23756; ROM4[6944]<=16'd57267;
ROM1[6945]<=16'd4750; ROM2[6945]<=16'd0; ROM3[6945]<=16'd23762; ROM4[6945]<=16'd57265;
ROM1[6946]<=16'd4750; ROM2[6946]<=16'd0; ROM3[6946]<=16'd23762; ROM4[6946]<=16'd57268;
ROM1[6947]<=16'd4793; ROM2[6947]<=16'd0; ROM3[6947]<=16'd23776; ROM4[6947]<=16'd57288;
ROM1[6948]<=16'd4861; ROM2[6948]<=16'd0; ROM3[6948]<=16'd23799; ROM4[6948]<=16'd57322;
ROM1[6949]<=16'd4863; ROM2[6949]<=16'd0; ROM3[6949]<=16'd23790; ROM4[6949]<=16'd57318;
ROM1[6950]<=16'd4809; ROM2[6950]<=16'd0; ROM3[6950]<=16'd23755; ROM4[6950]<=16'd57280;
ROM1[6951]<=16'd4763; ROM2[6951]<=16'd0; ROM3[6951]<=16'd23731; ROM4[6951]<=16'd57249;
ROM1[6952]<=16'd4739; ROM2[6952]<=16'd0; ROM3[6952]<=16'd23729; ROM4[6952]<=16'd57241;
ROM1[6953]<=16'd4726; ROM2[6953]<=16'd0; ROM3[6953]<=16'd23742; ROM4[6953]<=16'd57243;
ROM1[6954]<=16'd4738; ROM2[6954]<=16'd0; ROM3[6954]<=16'd23759; ROM4[6954]<=16'd57260;
ROM1[6955]<=16'd4758; ROM2[6955]<=16'd0; ROM3[6955]<=16'd23768; ROM4[6955]<=16'd57271;
ROM1[6956]<=16'd4778; ROM2[6956]<=16'd0; ROM3[6956]<=16'd23745; ROM4[6956]<=16'd57255;
ROM1[6957]<=16'd4801; ROM2[6957]<=16'd0; ROM3[6957]<=16'd23732; ROM4[6957]<=16'd57256;
ROM1[6958]<=16'd4814; ROM2[6958]<=16'd0; ROM3[6958]<=16'd23755; ROM4[6958]<=16'd57274;
ROM1[6959]<=16'd4800; ROM2[6959]<=16'd0; ROM3[6959]<=16'd23767; ROM4[6959]<=16'd57280;
ROM1[6960]<=16'd4769; ROM2[6960]<=16'd0; ROM3[6960]<=16'd23757; ROM4[6960]<=16'd57268;
ROM1[6961]<=16'd4749; ROM2[6961]<=16'd0; ROM3[6961]<=16'd23760; ROM4[6961]<=16'd57258;
ROM1[6962]<=16'd4725; ROM2[6962]<=16'd0; ROM3[6962]<=16'd23754; ROM4[6962]<=16'd57246;
ROM1[6963]<=16'd4729; ROM2[6963]<=16'd0; ROM3[6963]<=16'd23743; ROM4[6963]<=16'd57240;
ROM1[6964]<=16'd4764; ROM2[6964]<=16'd0; ROM3[6964]<=16'd23741; ROM4[6964]<=16'd57246;
ROM1[6965]<=16'd4798; ROM2[6965]<=16'd0; ROM3[6965]<=16'd23727; ROM4[6965]<=16'd57247;
ROM1[6966]<=16'd4799; ROM2[6966]<=16'd0; ROM3[6966]<=16'd23722; ROM4[6966]<=16'd57241;
ROM1[6967]<=16'd4778; ROM2[6967]<=16'd0; ROM3[6967]<=16'd23723; ROM4[6967]<=16'd57238;
ROM1[6968]<=16'd4759; ROM2[6968]<=16'd0; ROM3[6968]<=16'd23734; ROM4[6968]<=16'd57240;
ROM1[6969]<=16'd4741; ROM2[6969]<=16'd0; ROM3[6969]<=16'd23743; ROM4[6969]<=16'd57244;
ROM1[6970]<=16'd4728; ROM2[6970]<=16'd0; ROM3[6970]<=16'd23751; ROM4[6970]<=16'd57245;
ROM1[6971]<=16'd4730; ROM2[6971]<=16'd0; ROM3[6971]<=16'd23757; ROM4[6971]<=16'd57244;
ROM1[6972]<=16'd4751; ROM2[6972]<=16'd0; ROM3[6972]<=16'd23753; ROM4[6972]<=16'd57240;
ROM1[6973]<=16'd4786; ROM2[6973]<=16'd0; ROM3[6973]<=16'd23738; ROM4[6973]<=16'd57240;
ROM1[6974]<=16'd4798; ROM2[6974]<=16'd0; ROM3[6974]<=16'd23731; ROM4[6974]<=16'd57242;
ROM1[6975]<=16'd4787; ROM2[6975]<=16'd0; ROM3[6975]<=16'd23744; ROM4[6975]<=16'd57248;
ROM1[6976]<=16'd4769; ROM2[6976]<=16'd0; ROM3[6976]<=16'd23753; ROM4[6976]<=16'd57252;
ROM1[6977]<=16'd4758; ROM2[6977]<=16'd0; ROM3[6977]<=16'd23761; ROM4[6977]<=16'd57251;
ROM1[6978]<=16'd4748; ROM2[6978]<=16'd0; ROM3[6978]<=16'd23775; ROM4[6978]<=16'd57256;
ROM1[6979]<=16'd4731; ROM2[6979]<=16'd0; ROM3[6979]<=16'd23766; ROM4[6979]<=16'd57247;
ROM1[6980]<=16'd4749; ROM2[6980]<=16'd0; ROM3[6980]<=16'd23762; ROM4[6980]<=16'd57249;
ROM1[6981]<=16'd4787; ROM2[6981]<=16'd0; ROM3[6981]<=16'd23763; ROM4[6981]<=16'd57265;
ROM1[6982]<=16'd4806; ROM2[6982]<=16'd0; ROM3[6982]<=16'd23755; ROM4[6982]<=16'd57269;
ROM1[6983]<=16'd4793; ROM2[6983]<=16'd0; ROM3[6983]<=16'd23751; ROM4[6983]<=16'd57263;
ROM1[6984]<=16'd4772; ROM2[6984]<=16'd0; ROM3[6984]<=16'd23753; ROM4[6984]<=16'd57257;
ROM1[6985]<=16'd4762; ROM2[6985]<=16'd0; ROM3[6985]<=16'd23759; ROM4[6985]<=16'd57258;
ROM1[6986]<=16'd4746; ROM2[6986]<=16'd0; ROM3[6986]<=16'd23760; ROM4[6986]<=16'd57255;
ROM1[6987]<=16'd4735; ROM2[6987]<=16'd0; ROM3[6987]<=16'd23763; ROM4[6987]<=16'd57254;
ROM1[6988]<=16'd4740; ROM2[6988]<=16'd0; ROM3[6988]<=16'd23756; ROM4[6988]<=16'd57252;
ROM1[6989]<=16'd4753; ROM2[6989]<=16'd0; ROM3[6989]<=16'd23738; ROM4[6989]<=16'd57242;
ROM1[6990]<=16'd4784; ROM2[6990]<=16'd0; ROM3[6990]<=16'd23733; ROM4[6990]<=16'd57244;
ROM1[6991]<=16'd4800; ROM2[6991]<=16'd0; ROM3[6991]<=16'd23743; ROM4[6991]<=16'd57257;
ROM1[6992]<=16'd4791; ROM2[6992]<=16'd0; ROM3[6992]<=16'd23755; ROM4[6992]<=16'd57264;
ROM1[6993]<=16'd4774; ROM2[6993]<=16'd0; ROM3[6993]<=16'd23769; ROM4[6993]<=16'd57262;
ROM1[6994]<=16'd4766; ROM2[6994]<=16'd0; ROM3[6994]<=16'd23778; ROM4[6994]<=16'd57270;
ROM1[6995]<=16'd4766; ROM2[6995]<=16'd0; ROM3[6995]<=16'd23795; ROM4[6995]<=16'd57283;
ROM1[6996]<=16'd4759; ROM2[6996]<=16'd0; ROM3[6996]<=16'd23786; ROM4[6996]<=16'd57276;
ROM1[6997]<=16'd4767; ROM2[6997]<=16'd0; ROM3[6997]<=16'd23762; ROM4[6997]<=16'd57265;
ROM1[6998]<=16'd4805; ROM2[6998]<=16'd0; ROM3[6998]<=16'd23756; ROM4[6998]<=16'd57267;
ROM1[6999]<=16'd4811; ROM2[6999]<=16'd0; ROM3[6999]<=16'd23747; ROM4[6999]<=16'd57262;
ROM1[7000]<=16'd4786; ROM2[7000]<=16'd0; ROM3[7000]<=16'd23744; ROM4[7000]<=16'd57254;
ROM1[7001]<=16'd4789; ROM2[7001]<=16'd0; ROM3[7001]<=16'd23772; ROM4[7001]<=16'd57275;
ROM1[7002]<=16'd4772; ROM2[7002]<=16'd0; ROM3[7002]<=16'd23771; ROM4[7002]<=16'd57267;
ROM1[7003]<=16'd4734; ROM2[7003]<=16'd0; ROM3[7003]<=16'd23750; ROM4[7003]<=16'd57240;
ROM1[7004]<=16'd4730; ROM2[7004]<=16'd0; ROM3[7004]<=16'd23753; ROM4[7004]<=16'd57242;
ROM1[7005]<=16'd4753; ROM2[7005]<=16'd0; ROM3[7005]<=16'd23758; ROM4[7005]<=16'd57250;
ROM1[7006]<=16'd4805; ROM2[7006]<=16'd0; ROM3[7006]<=16'd23763; ROM4[7006]<=16'd57267;
ROM1[7007]<=16'd4836; ROM2[7007]<=16'd0; ROM3[7007]<=16'd23760; ROM4[7007]<=16'd57276;
ROM1[7008]<=16'd4817; ROM2[7008]<=16'd0; ROM3[7008]<=16'd23753; ROM4[7008]<=16'd57263;
ROM1[7009]<=16'd4779; ROM2[7009]<=16'd0; ROM3[7009]<=16'd23742; ROM4[7009]<=16'd57244;
ROM1[7010]<=16'd4752; ROM2[7010]<=16'd0; ROM3[7010]<=16'd23742; ROM4[7010]<=16'd57238;
ROM1[7011]<=16'd4747; ROM2[7011]<=16'd0; ROM3[7011]<=16'd23758; ROM4[7011]<=16'd57243;
ROM1[7012]<=16'd4752; ROM2[7012]<=16'd0; ROM3[7012]<=16'd23774; ROM4[7012]<=16'd57258;
ROM1[7013]<=16'd4764; ROM2[7013]<=16'd0; ROM3[7013]<=16'd23777; ROM4[7013]<=16'd57266;
ROM1[7014]<=16'd4787; ROM2[7014]<=16'd0; ROM3[7014]<=16'd23765; ROM4[7014]<=16'd57260;
ROM1[7015]<=16'd4816; ROM2[7015]<=16'd0; ROM3[7015]<=16'd23758; ROM4[7015]<=16'd57261;
ROM1[7016]<=16'd4821; ROM2[7016]<=16'd0; ROM3[7016]<=16'd23762; ROM4[7016]<=16'd57267;
ROM1[7017]<=16'd4804; ROM2[7017]<=16'd0; ROM3[7017]<=16'd23766; ROM4[7017]<=16'd57266;
ROM1[7018]<=16'd4781; ROM2[7018]<=16'd0; ROM3[7018]<=16'd23767; ROM4[7018]<=16'd57263;
ROM1[7019]<=16'd4764; ROM2[7019]<=16'd0; ROM3[7019]<=16'd23767; ROM4[7019]<=16'd57264;
ROM1[7020]<=16'd4754; ROM2[7020]<=16'd0; ROM3[7020]<=16'd23779; ROM4[7020]<=16'd57269;
ROM1[7021]<=16'd4757; ROM2[7021]<=16'd0; ROM3[7021]<=16'd23776; ROM4[7021]<=16'd57269;
ROM1[7022]<=16'd4781; ROM2[7022]<=16'd0; ROM3[7022]<=16'd23766; ROM4[7022]<=16'd57268;
ROM1[7023]<=16'd4810; ROM2[7023]<=16'd0; ROM3[7023]<=16'd23745; ROM4[7023]<=16'd57263;
ROM1[7024]<=16'd4815; ROM2[7024]<=16'd0; ROM3[7024]<=16'd23733; ROM4[7024]<=16'd57256;
ROM1[7025]<=16'd4802; ROM2[7025]<=16'd0; ROM3[7025]<=16'd23735; ROM4[7025]<=16'd57252;
ROM1[7026]<=16'd4790; ROM2[7026]<=16'd0; ROM3[7026]<=16'd23748; ROM4[7026]<=16'd57258;
ROM1[7027]<=16'd4790; ROM2[7027]<=16'd0; ROM3[7027]<=16'd23771; ROM4[7027]<=16'd57273;
ROM1[7028]<=16'd4781; ROM2[7028]<=16'd0; ROM3[7028]<=16'd23781; ROM4[7028]<=16'd57277;
ROM1[7029]<=16'd4768; ROM2[7029]<=16'd0; ROM3[7029]<=16'd23779; ROM4[7029]<=16'd57275;
ROM1[7030]<=16'd4780; ROM2[7030]<=16'd0; ROM3[7030]<=16'd23778; ROM4[7030]<=16'd57274;
ROM1[7031]<=16'd4816; ROM2[7031]<=16'd0; ROM3[7031]<=16'd23770; ROM4[7031]<=16'd57274;
ROM1[7032]<=16'd4838; ROM2[7032]<=16'd0; ROM3[7032]<=16'd23764; ROM4[7032]<=16'd57273;
ROM1[7033]<=16'd4835; ROM2[7033]<=16'd0; ROM3[7033]<=16'd23778; ROM4[7033]<=16'd57281;
ROM1[7034]<=16'd4812; ROM2[7034]<=16'd0; ROM3[7034]<=16'd23784; ROM4[7034]<=16'd57279;
ROM1[7035]<=16'd4784; ROM2[7035]<=16'd0; ROM3[7035]<=16'd23779; ROM4[7035]<=16'd57264;
ROM1[7036]<=16'd4769; ROM2[7036]<=16'd0; ROM3[7036]<=16'd23782; ROM4[7036]<=16'd57265;
ROM1[7037]<=16'd4769; ROM2[7037]<=16'd0; ROM3[7037]<=16'd23796; ROM4[7037]<=16'd57276;
ROM1[7038]<=16'd4791; ROM2[7038]<=16'd0; ROM3[7038]<=16'd23808; ROM4[7038]<=16'd57290;
ROM1[7039]<=16'd4819; ROM2[7039]<=16'd0; ROM3[7039]<=16'd23797; ROM4[7039]<=16'd57292;
ROM1[7040]<=16'd4846; ROM2[7040]<=16'd0; ROM3[7040]<=16'd23783; ROM4[7040]<=16'd57288;
ROM1[7041]<=16'd4822; ROM2[7041]<=16'd0; ROM3[7041]<=16'd23753; ROM4[7041]<=16'd57265;
ROM1[7042]<=16'd4797; ROM2[7042]<=16'd0; ROM3[7042]<=16'd23749; ROM4[7042]<=16'd57261;
ROM1[7043]<=16'd4788; ROM2[7043]<=16'd0; ROM3[7043]<=16'd23766; ROM4[7043]<=16'd57273;
ROM1[7044]<=16'd4781; ROM2[7044]<=16'd0; ROM3[7044]<=16'd23777; ROM4[7044]<=16'd57280;
ROM1[7045]<=16'd4787; ROM2[7045]<=16'd0; ROM3[7045]<=16'd23796; ROM4[7045]<=16'd57294;
ROM1[7046]<=16'd4782; ROM2[7046]<=16'd0; ROM3[7046]<=16'd23791; ROM4[7046]<=16'd57284;
ROM1[7047]<=16'd4787; ROM2[7047]<=16'd0; ROM3[7047]<=16'd23772; ROM4[7047]<=16'd57272;
ROM1[7048]<=16'd4813; ROM2[7048]<=16'd0; ROM3[7048]<=16'd23758; ROM4[7048]<=16'd57269;
ROM1[7049]<=16'd4825; ROM2[7049]<=16'd0; ROM3[7049]<=16'd23751; ROM4[7049]<=16'd57267;
ROM1[7050]<=16'd4817; ROM2[7050]<=16'd0; ROM3[7050]<=16'd23758; ROM4[7050]<=16'd57271;
ROM1[7051]<=16'd4805; ROM2[7051]<=16'd0; ROM3[7051]<=16'd23770; ROM4[7051]<=16'd57276;
ROM1[7052]<=16'd4794; ROM2[7052]<=16'd0; ROM3[7052]<=16'd23777; ROM4[7052]<=16'd57278;
ROM1[7053]<=16'd4777; ROM2[7053]<=16'd0; ROM3[7053]<=16'd23786; ROM4[7053]<=16'd57278;
ROM1[7054]<=16'd4769; ROM2[7054]<=16'd0; ROM3[7054]<=16'd23784; ROM4[7054]<=16'd57277;
ROM1[7055]<=16'd4784; ROM2[7055]<=16'd0; ROM3[7055]<=16'd23776; ROM4[7055]<=16'd57274;
ROM1[7056]<=16'd4819; ROM2[7056]<=16'd0; ROM3[7056]<=16'd23764; ROM4[7056]<=16'd57273;
ROM1[7057]<=16'd4843; ROM2[7057]<=16'd0; ROM3[7057]<=16'd23761; ROM4[7057]<=16'd57274;
ROM1[7058]<=16'd4837; ROM2[7058]<=16'd0; ROM3[7058]<=16'd23772; ROM4[7058]<=16'd57280;
ROM1[7059]<=16'd4816; ROM2[7059]<=16'd0; ROM3[7059]<=16'd23780; ROM4[7059]<=16'd57278;
ROM1[7060]<=16'd4800; ROM2[7060]<=16'd0; ROM3[7060]<=16'd23794; ROM4[7060]<=16'd57280;
ROM1[7061]<=16'd4793; ROM2[7061]<=16'd0; ROM3[7061]<=16'd23810; ROM4[7061]<=16'd57289;
ROM1[7062]<=16'd4766; ROM2[7062]<=16'd0; ROM3[7062]<=16'd23801; ROM4[7062]<=16'd57277;
ROM1[7063]<=16'd4765; ROM2[7063]<=16'd0; ROM3[7063]<=16'd23797; ROM4[7063]<=16'd57274;
ROM1[7064]<=16'd4797; ROM2[7064]<=16'd0; ROM3[7064]<=16'd23782; ROM4[7064]<=16'd57271;
ROM1[7065]<=16'd4831; ROM2[7065]<=16'd0; ROM3[7065]<=16'd23761; ROM4[7065]<=16'd57265;
ROM1[7066]<=16'd4844; ROM2[7066]<=16'd0; ROM3[7066]<=16'd23768; ROM4[7066]<=16'd57272;
ROM1[7067]<=16'd4828; ROM2[7067]<=16'd0; ROM3[7067]<=16'd23773; ROM4[7067]<=16'd57277;
ROM1[7068]<=16'd4808; ROM2[7068]<=16'd0; ROM3[7068]<=16'd23779; ROM4[7068]<=16'd57278;
ROM1[7069]<=16'd4790; ROM2[7069]<=16'd0; ROM3[7069]<=16'd23780; ROM4[7069]<=16'd57273;
ROM1[7070]<=16'd4775; ROM2[7070]<=16'd0; ROM3[7070]<=16'd23777; ROM4[7070]<=16'd57267;
ROM1[7071]<=16'd4781; ROM2[7071]<=16'd0; ROM3[7071]<=16'd23779; ROM4[7071]<=16'd57264;
ROM1[7072]<=16'd4801; ROM2[7072]<=16'd0; ROM3[7072]<=16'd23776; ROM4[7072]<=16'd57267;
ROM1[7073]<=16'd4830; ROM2[7073]<=16'd0; ROM3[7073]<=16'd23765; ROM4[7073]<=16'd57272;
ROM1[7074]<=16'd4858; ROM2[7074]<=16'd0; ROM3[7074]<=16'd23780; ROM4[7074]<=16'd57295;
ROM1[7075]<=16'd4855; ROM2[7075]<=16'd0; ROM3[7075]<=16'd23793; ROM4[7075]<=16'd57305;
ROM1[7076]<=16'd4812; ROM2[7076]<=16'd0; ROM3[7076]<=16'd23780; ROM4[7076]<=16'd57285;
ROM1[7077]<=16'd4782; ROM2[7077]<=16'd0; ROM3[7077]<=16'd23776; ROM4[7077]<=16'd57273;
ROM1[7078]<=16'd4768; ROM2[7078]<=16'd0; ROM3[7078]<=16'd23780; ROM4[7078]<=16'd57270;
ROM1[7079]<=16'd4767; ROM2[7079]<=16'd0; ROM3[7079]<=16'd23791; ROM4[7079]<=16'd57277;
ROM1[7080]<=16'd4795; ROM2[7080]<=16'd0; ROM3[7080]<=16'd23806; ROM4[7080]<=16'd57294;
ROM1[7081]<=16'd4824; ROM2[7081]<=16'd0; ROM3[7081]<=16'd23794; ROM4[7081]<=16'd57290;
ROM1[7082]<=16'd4831; ROM2[7082]<=16'd0; ROM3[7082]<=16'd23770; ROM4[7082]<=16'd57273;
ROM1[7083]<=16'd4812; ROM2[7083]<=16'd0; ROM3[7083]<=16'd23757; ROM4[7083]<=16'd57263;
ROM1[7084]<=16'd4789; ROM2[7084]<=16'd0; ROM3[7084]<=16'd23759; ROM4[7084]<=16'd57259;
ROM1[7085]<=16'd4782; ROM2[7085]<=16'd0; ROM3[7085]<=16'd23774; ROM4[7085]<=16'd57261;
ROM1[7086]<=16'd4776; ROM2[7086]<=16'd0; ROM3[7086]<=16'd23786; ROM4[7086]<=16'd57269;
ROM1[7087]<=16'd4787; ROM2[7087]<=16'd0; ROM3[7087]<=16'd23804; ROM4[7087]<=16'd57287;
ROM1[7088]<=16'd4808; ROM2[7088]<=16'd0; ROM3[7088]<=16'd23812; ROM4[7088]<=16'd57297;
ROM1[7089]<=16'd4815; ROM2[7089]<=16'd0; ROM3[7089]<=16'd23781; ROM4[7089]<=16'd57276;
ROM1[7090]<=16'd4821; ROM2[7090]<=16'd0; ROM3[7090]<=16'd23748; ROM4[7090]<=16'd57250;
ROM1[7091]<=16'd4812; ROM2[7091]<=16'd0; ROM3[7091]<=16'd23740; ROM4[7091]<=16'd57243;
ROM1[7092]<=16'd4795; ROM2[7092]<=16'd0; ROM3[7092]<=16'd23744; ROM4[7092]<=16'd57246;
ROM1[7093]<=16'd4780; ROM2[7093]<=16'd0; ROM3[7093]<=16'd23753; ROM4[7093]<=16'd57253;
ROM1[7094]<=16'd4762; ROM2[7094]<=16'd0; ROM3[7094]<=16'd23756; ROM4[7094]<=16'd57254;
ROM1[7095]<=16'd4738; ROM2[7095]<=16'd0; ROM3[7095]<=16'd23749; ROM4[7095]<=16'd57244;
ROM1[7096]<=16'd4733; ROM2[7096]<=16'd0; ROM3[7096]<=16'd23742; ROM4[7096]<=16'd57239;
ROM1[7097]<=16'd4762; ROM2[7097]<=16'd0; ROM3[7097]<=16'd23742; ROM4[7097]<=16'd57248;
ROM1[7098]<=16'd4802; ROM2[7098]<=16'd0; ROM3[7098]<=16'd23740; ROM4[7098]<=16'd57258;
ROM1[7099]<=16'd4817; ROM2[7099]<=16'd0; ROM3[7099]<=16'd23742; ROM4[7099]<=16'd57263;
ROM1[7100]<=16'd4802; ROM2[7100]<=16'd0; ROM3[7100]<=16'd23746; ROM4[7100]<=16'd57259;
ROM1[7101]<=16'd4794; ROM2[7101]<=16'd0; ROM3[7101]<=16'd23759; ROM4[7101]<=16'd57262;
ROM1[7102]<=16'd4789; ROM2[7102]<=16'd0; ROM3[7102]<=16'd23775; ROM4[7102]<=16'd57275;
ROM1[7103]<=16'd4778; ROM2[7103]<=16'd0; ROM3[7103]<=16'd23781; ROM4[7103]<=16'd57275;
ROM1[7104]<=16'd4779; ROM2[7104]<=16'd0; ROM3[7104]<=16'd23789; ROM4[7104]<=16'd57281;
ROM1[7105]<=16'd4786; ROM2[7105]<=16'd0; ROM3[7105]<=16'd23785; ROM4[7105]<=16'd57279;
ROM1[7106]<=16'd4809; ROM2[7106]<=16'd0; ROM3[7106]<=16'd23772; ROM4[7106]<=16'd57268;
ROM1[7107]<=16'd4821; ROM2[7107]<=16'd0; ROM3[7107]<=16'd23760; ROM4[7107]<=16'd57265;
ROM1[7108]<=16'd4811; ROM2[7108]<=16'd0; ROM3[7108]<=16'd23762; ROM4[7108]<=16'd57267;
ROM1[7109]<=16'd4809; ROM2[7109]<=16'd0; ROM3[7109]<=16'd23781; ROM4[7109]<=16'd57279;
ROM1[7110]<=16'd4798; ROM2[7110]<=16'd0; ROM3[7110]<=16'd23788; ROM4[7110]<=16'd57281;
ROM1[7111]<=16'd4783; ROM2[7111]<=16'd0; ROM3[7111]<=16'd23792; ROM4[7111]<=16'd57279;
ROM1[7112]<=16'd4776; ROM2[7112]<=16'd0; ROM3[7112]<=16'd23796; ROM4[7112]<=16'd57283;
ROM1[7113]<=16'd4781; ROM2[7113]<=16'd0; ROM3[7113]<=16'd23795; ROM4[7113]<=16'd57288;
ROM1[7114]<=16'd4816; ROM2[7114]<=16'd0; ROM3[7114]<=16'd23794; ROM4[7114]<=16'd57295;
ROM1[7115]<=16'd4849; ROM2[7115]<=16'd0; ROM3[7115]<=16'd23790; ROM4[7115]<=16'd57302;
ROM1[7116]<=16'd4840; ROM2[7116]<=16'd0; ROM3[7116]<=16'd23786; ROM4[7116]<=16'd57294;
ROM1[7117]<=16'd4819; ROM2[7117]<=16'd0; ROM3[7117]<=16'd23781; ROM4[7117]<=16'd57284;
ROM1[7118]<=16'd4801; ROM2[7118]<=16'd0; ROM3[7118]<=16'd23790; ROM4[7118]<=16'd57289;
ROM1[7119]<=16'd4794; ROM2[7119]<=16'd0; ROM3[7119]<=16'd23802; ROM4[7119]<=16'd57295;
ROM1[7120]<=16'd4777; ROM2[7120]<=16'd0; ROM3[7120]<=16'd23797; ROM4[7120]<=16'd57286;
ROM1[7121]<=16'd4774; ROM2[7121]<=16'd0; ROM3[7121]<=16'd23793; ROM4[7121]<=16'd57278;
ROM1[7122]<=16'd4793; ROM2[7122]<=16'd0; ROM3[7122]<=16'd23784; ROM4[7122]<=16'd57275;
ROM1[7123]<=16'd4821; ROM2[7123]<=16'd0; ROM3[7123]<=16'd23770; ROM4[7123]<=16'd57271;
ROM1[7124]<=16'd4835; ROM2[7124]<=16'd0; ROM3[7124]<=16'd23772; ROM4[7124]<=16'd57277;
ROM1[7125]<=16'd4821; ROM2[7125]<=16'd0; ROM3[7125]<=16'd23775; ROM4[7125]<=16'd57278;
ROM1[7126]<=16'd4800; ROM2[7126]<=16'd0; ROM3[7126]<=16'd23776; ROM4[7126]<=16'd57275;
ROM1[7127]<=16'd4809; ROM2[7127]<=16'd0; ROM3[7127]<=16'd23797; ROM4[7127]<=16'd57295;
ROM1[7128]<=16'd4808; ROM2[7128]<=16'd0; ROM3[7128]<=16'd23815; ROM4[7128]<=16'd57311;
ROM1[7129]<=16'd4803; ROM2[7129]<=16'd0; ROM3[7129]<=16'd23819; ROM4[7129]<=16'd57315;
ROM1[7130]<=16'd4804; ROM2[7130]<=16'd0; ROM3[7130]<=16'd23805; ROM4[7130]<=16'd57304;
ROM1[7131]<=16'd4815; ROM2[7131]<=16'd0; ROM3[7131]<=16'd23770; ROM4[7131]<=16'd57280;
ROM1[7132]<=16'd4844; ROM2[7132]<=16'd0; ROM3[7132]<=16'd23761; ROM4[7132]<=16'd57281;
ROM1[7133]<=16'd4843; ROM2[7133]<=16'd0; ROM3[7133]<=16'd23766; ROM4[7133]<=16'd57284;
ROM1[7134]<=16'd4823; ROM2[7134]<=16'd0; ROM3[7134]<=16'd23770; ROM4[7134]<=16'd57284;
ROM1[7135]<=16'd4808; ROM2[7135]<=16'd0; ROM3[7135]<=16'd23782; ROM4[7135]<=16'd57289;
ROM1[7136]<=16'd4788; ROM2[7136]<=16'd0; ROM3[7136]<=16'd23779; ROM4[7136]<=16'd57281;
ROM1[7137]<=16'd4777; ROM2[7137]<=16'd0; ROM3[7137]<=16'd23779; ROM4[7137]<=16'd57274;
ROM1[7138]<=16'd4789; ROM2[7138]<=16'd0; ROM3[7138]<=16'd23777; ROM4[7138]<=16'd57276;
ROM1[7139]<=16'd4819; ROM2[7139]<=16'd0; ROM3[7139]<=16'd23766; ROM4[7139]<=16'd57279;
ROM1[7140]<=16'd4838; ROM2[7140]<=16'd0; ROM3[7140]<=16'd23756; ROM4[7140]<=16'd57274;
ROM1[7141]<=16'd4820; ROM2[7141]<=16'd0; ROM3[7141]<=16'd23739; ROM4[7141]<=16'd57259;
ROM1[7142]<=16'd4801; ROM2[7142]<=16'd0; ROM3[7142]<=16'd23744; ROM4[7142]<=16'd57256;
ROM1[7143]<=16'd4775; ROM2[7143]<=16'd0; ROM3[7143]<=16'd23748; ROM4[7143]<=16'd57250;
ROM1[7144]<=16'd4756; ROM2[7144]<=16'd0; ROM3[7144]<=16'd23750; ROM4[7144]<=16'd57248;
ROM1[7145]<=16'd4758; ROM2[7145]<=16'd0; ROM3[7145]<=16'd23768; ROM4[7145]<=16'd57261;
ROM1[7146]<=16'd4764; ROM2[7146]<=16'd0; ROM3[7146]<=16'd23770; ROM4[7146]<=16'd57260;
ROM1[7147]<=16'd4781; ROM2[7147]<=16'd0; ROM3[7147]<=16'd23756; ROM4[7147]<=16'd57252;
ROM1[7148]<=16'd4805; ROM2[7148]<=16'd0; ROM3[7148]<=16'd23738; ROM4[7148]<=16'd57240;
ROM1[7149]<=16'd4818; ROM2[7149]<=16'd0; ROM3[7149]<=16'd23742; ROM4[7149]<=16'd57250;
ROM1[7150]<=16'd4809; ROM2[7150]<=16'd0; ROM3[7150]<=16'd23754; ROM4[7150]<=16'd57259;
ROM1[7151]<=16'd4796; ROM2[7151]<=16'd0; ROM3[7151]<=16'd23772; ROM4[7151]<=16'd57264;
ROM1[7152]<=16'd4800; ROM2[7152]<=16'd0; ROM3[7152]<=16'd23794; ROM4[7152]<=16'd57283;
ROM1[7153]<=16'd4798; ROM2[7153]<=16'd0; ROM3[7153]<=16'd23804; ROM4[7153]<=16'd57286;
ROM1[7154]<=16'd4780; ROM2[7154]<=16'd0; ROM3[7154]<=16'd23785; ROM4[7154]<=16'd57267;
ROM1[7155]<=16'd4781; ROM2[7155]<=16'd0; ROM3[7155]<=16'd23765; ROM4[7155]<=16'd57253;
ROM1[7156]<=16'd4811; ROM2[7156]<=16'd0; ROM3[7156]<=16'd23757; ROM4[7156]<=16'd57255;
ROM1[7157]<=16'd4819; ROM2[7157]<=16'd0; ROM3[7157]<=16'd23739; ROM4[7157]<=16'd57249;
ROM1[7158]<=16'd4810; ROM2[7158]<=16'd0; ROM3[7158]<=16'd23746; ROM4[7158]<=16'd57251;
ROM1[7159]<=16'd4799; ROM2[7159]<=16'd0; ROM3[7159]<=16'd23757; ROM4[7159]<=16'd57254;
ROM1[7160]<=16'd4782; ROM2[7160]<=16'd0; ROM3[7160]<=16'd23755; ROM4[7160]<=16'd57247;
ROM1[7161]<=16'd4772; ROM2[7161]<=16'd0; ROM3[7161]<=16'd23771; ROM4[7161]<=16'd57253;
ROM1[7162]<=16'd4767; ROM2[7162]<=16'd0; ROM3[7162]<=16'd23778; ROM4[7162]<=16'd57261;
ROM1[7163]<=16'd4775; ROM2[7163]<=16'd0; ROM3[7163]<=16'd23774; ROM4[7163]<=16'd57263;
ROM1[7164]<=16'd4798; ROM2[7164]<=16'd0; ROM3[7164]<=16'd23765; ROM4[7164]<=16'd57262;
ROM1[7165]<=16'd4825; ROM2[7165]<=16'd0; ROM3[7165]<=16'd23753; ROM4[7165]<=16'd57263;
ROM1[7166]<=16'd4834; ROM2[7166]<=16'd0; ROM3[7166]<=16'd23765; ROM4[7166]<=16'd57271;
ROM1[7167]<=16'd4824; ROM2[7167]<=16'd0; ROM3[7167]<=16'd23781; ROM4[7167]<=16'd57281;
ROM1[7168]<=16'd4804; ROM2[7168]<=16'd0; ROM3[7168]<=16'd23791; ROM4[7168]<=16'd57286;
ROM1[7169]<=16'd4787; ROM2[7169]<=16'd0; ROM3[7169]<=16'd23797; ROM4[7169]<=16'd57284;
ROM1[7170]<=16'd4766; ROM2[7170]<=16'd0; ROM3[7170]<=16'd23793; ROM4[7170]<=16'd57276;
ROM1[7171]<=16'd4759; ROM2[7171]<=16'd0; ROM3[7171]<=16'd23784; ROM4[7171]<=16'd57267;
ROM1[7172]<=16'd4778; ROM2[7172]<=16'd0; ROM3[7172]<=16'd23774; ROM4[7172]<=16'd57262;
ROM1[7173]<=16'd4803; ROM2[7173]<=16'd0; ROM3[7173]<=16'd23759; ROM4[7173]<=16'd57260;
ROM1[7174]<=16'd4804; ROM2[7174]<=16'd0; ROM3[7174]<=16'd23750; ROM4[7174]<=16'd57253;
ROM1[7175]<=16'd4790; ROM2[7175]<=16'd0; ROM3[7175]<=16'd23756; ROM4[7175]<=16'd57251;
ROM1[7176]<=16'd4778; ROM2[7176]<=16'd0; ROM3[7176]<=16'd23765; ROM4[7176]<=16'd57254;
ROM1[7177]<=16'd4766; ROM2[7177]<=16'd0; ROM3[7177]<=16'd23771; ROM4[7177]<=16'd57254;
ROM1[7178]<=16'd4752; ROM2[7178]<=16'd0; ROM3[7178]<=16'd23782; ROM4[7178]<=16'd57260;
ROM1[7179]<=16'd4754; ROM2[7179]<=16'd0; ROM3[7179]<=16'd23791; ROM4[7179]<=16'd57268;
ROM1[7180]<=16'd4768; ROM2[7180]<=16'd0; ROM3[7180]<=16'd23787; ROM4[7180]<=16'd57266;
ROM1[7181]<=16'd4800; ROM2[7181]<=16'd0; ROM3[7181]<=16'd23775; ROM4[7181]<=16'd57265;
ROM1[7182]<=16'd4826; ROM2[7182]<=16'd0; ROM3[7182]<=16'd23767; ROM4[7182]<=16'd57262;
ROM1[7183]<=16'd4810; ROM2[7183]<=16'd0; ROM3[7183]<=16'd23764; ROM4[7183]<=16'd57255;
ROM1[7184]<=16'd4785; ROM2[7184]<=16'd0; ROM3[7184]<=16'd23768; ROM4[7184]<=16'd57253;
ROM1[7185]<=16'd4771; ROM2[7185]<=16'd0; ROM3[7185]<=16'd23779; ROM4[7185]<=16'd57254;
ROM1[7186]<=16'd4772; ROM2[7186]<=16'd0; ROM3[7186]<=16'd23795; ROM4[7186]<=16'd57272;
ROM1[7187]<=16'd4777; ROM2[7187]<=16'd0; ROM3[7187]<=16'd23806; ROM4[7187]<=16'd57284;
ROM1[7188]<=16'd4776; ROM2[7188]<=16'd0; ROM3[7188]<=16'd23793; ROM4[7188]<=16'd57275;
ROM1[7189]<=16'd4785; ROM2[7189]<=16'd0; ROM3[7189]<=16'd23767; ROM4[7189]<=16'd57261;
ROM1[7190]<=16'd4807; ROM2[7190]<=16'd0; ROM3[7190]<=16'd23755; ROM4[7190]<=16'd57258;
ROM1[7191]<=16'd4806; ROM2[7191]<=16'd0; ROM3[7191]<=16'd23757; ROM4[7191]<=16'd57260;
ROM1[7192]<=16'd4786; ROM2[7192]<=16'd0; ROM3[7192]<=16'd23760; ROM4[7192]<=16'd57257;
ROM1[7193]<=16'd4779; ROM2[7193]<=16'd0; ROM3[7193]<=16'd23779; ROM4[7193]<=16'd57266;
ROM1[7194]<=16'd4785; ROM2[7194]<=16'd0; ROM3[7194]<=16'd23802; ROM4[7194]<=16'd57286;
ROM1[7195]<=16'd4772; ROM2[7195]<=16'd0; ROM3[7195]<=16'd23805; ROM4[7195]<=16'd57283;
ROM1[7196]<=16'd4767; ROM2[7196]<=16'd0; ROM3[7196]<=16'd23796; ROM4[7196]<=16'd57277;
ROM1[7197]<=16'd4783; ROM2[7197]<=16'd0; ROM3[7197]<=16'd23784; ROM4[7197]<=16'd57272;
ROM1[7198]<=16'd4794; ROM2[7198]<=16'd0; ROM3[7198]<=16'd23755; ROM4[7198]<=16'd57252;
ROM1[7199]<=16'd4806; ROM2[7199]<=16'd0; ROM3[7199]<=16'd23754; ROM4[7199]<=16'd57255;
ROM1[7200]<=16'd4806; ROM2[7200]<=16'd0; ROM3[7200]<=16'd23765; ROM4[7200]<=16'd57257;
ROM1[7201]<=16'd4784; ROM2[7201]<=16'd0; ROM3[7201]<=16'd23768; ROM4[7201]<=16'd57257;
ROM1[7202]<=16'd4778; ROM2[7202]<=16'd0; ROM3[7202]<=16'd23783; ROM4[7202]<=16'd57267;
ROM1[7203]<=16'd4762; ROM2[7203]<=16'd0; ROM3[7203]<=16'd23786; ROM4[7203]<=16'd57261;
ROM1[7204]<=16'd4763; ROM2[7204]<=16'd0; ROM3[7204]<=16'd23795; ROM4[7204]<=16'd57270;
ROM1[7205]<=16'd4794; ROM2[7205]<=16'd0; ROM3[7205]<=16'd23797; ROM4[7205]<=16'd57276;
ROM1[7206]<=16'd4820; ROM2[7206]<=16'd0; ROM3[7206]<=16'd23776; ROM4[7206]<=16'd57267;
ROM1[7207]<=16'd4828; ROM2[7207]<=16'd0; ROM3[7207]<=16'd23759; ROM4[7207]<=16'd57262;
ROM1[7208]<=16'd4811; ROM2[7208]<=16'd0; ROM3[7208]<=16'd23755; ROM4[7208]<=16'd57260;
ROM1[7209]<=16'd4792; ROM2[7209]<=16'd0; ROM3[7209]<=16'd23760; ROM4[7209]<=16'd57260;
ROM1[7210]<=16'd4773; ROM2[7210]<=16'd0; ROM3[7210]<=16'd23761; ROM4[7210]<=16'd57258;
ROM1[7211]<=16'd4764; ROM2[7211]<=16'd0; ROM3[7211]<=16'd23766; ROM4[7211]<=16'd57261;
ROM1[7212]<=16'd4770; ROM2[7212]<=16'd0; ROM3[7212]<=16'd23781; ROM4[7212]<=16'd57276;
ROM1[7213]<=16'd4775; ROM2[7213]<=16'd0; ROM3[7213]<=16'd23777; ROM4[7213]<=16'd57278;
ROM1[7214]<=16'd4792; ROM2[7214]<=16'd0; ROM3[7214]<=16'd23759; ROM4[7214]<=16'd57267;
ROM1[7215]<=16'd4826; ROM2[7215]<=16'd0; ROM3[7215]<=16'd23750; ROM4[7215]<=16'd57273;
ROM1[7216]<=16'd4829; ROM2[7216]<=16'd0; ROM3[7216]<=16'd23752; ROM4[7216]<=16'd57275;
ROM1[7217]<=16'd4812; ROM2[7217]<=16'd0; ROM3[7217]<=16'd23757; ROM4[7217]<=16'd57273;
ROM1[7218]<=16'd4796; ROM2[7218]<=16'd0; ROM3[7218]<=16'd23762; ROM4[7218]<=16'd57270;
ROM1[7219]<=16'd4783; ROM2[7219]<=16'd0; ROM3[7219]<=16'd23765; ROM4[7219]<=16'd57268;
ROM1[7220]<=16'd4785; ROM2[7220]<=16'd0; ROM3[7220]<=16'd23780; ROM4[7220]<=16'd57274;
ROM1[7221]<=16'd4809; ROM2[7221]<=16'd0; ROM3[7221]<=16'd23797; ROM4[7221]<=16'd57288;
ROM1[7222]<=16'd4838; ROM2[7222]<=16'd0; ROM3[7222]<=16'd23801; ROM4[7222]<=16'd57299;
ROM1[7223]<=16'd4853; ROM2[7223]<=16'd0; ROM3[7223]<=16'd23778; ROM4[7223]<=16'd57287;
ROM1[7224]<=16'd4843; ROM2[7224]<=16'd0; ROM3[7224]<=16'd23758; ROM4[7224]<=16'd57272;
ROM1[7225]<=16'd4821; ROM2[7225]<=16'd0; ROM3[7225]<=16'd23756; ROM4[7225]<=16'd57265;
ROM1[7226]<=16'd4806; ROM2[7226]<=16'd0; ROM3[7226]<=16'd23767; ROM4[7226]<=16'd57269;
ROM1[7227]<=16'd4804; ROM2[7227]<=16'd0; ROM3[7227]<=16'd23786; ROM4[7227]<=16'd57282;
ROM1[7228]<=16'd4775; ROM2[7228]<=16'd0; ROM3[7228]<=16'd23779; ROM4[7228]<=16'd57269;
ROM1[7229]<=16'd4762; ROM2[7229]<=16'd0; ROM3[7229]<=16'd23768; ROM4[7229]<=16'd57256;
ROM1[7230]<=16'd4772; ROM2[7230]<=16'd0; ROM3[7230]<=16'd23759; ROM4[7230]<=16'd57247;
ROM1[7231]<=16'd4791; ROM2[7231]<=16'd0; ROM3[7231]<=16'd23733; ROM4[7231]<=16'd57235;
ROM1[7232]<=16'd4819; ROM2[7232]<=16'd0; ROM3[7232]<=16'd23728; ROM4[7232]<=16'd57244;
ROM1[7233]<=16'd4818; ROM2[7233]<=16'd0; ROM3[7233]<=16'd23733; ROM4[7233]<=16'd57249;
ROM1[7234]<=16'd4808; ROM2[7234]<=16'd0; ROM3[7234]<=16'd23745; ROM4[7234]<=16'd57253;
ROM1[7235]<=16'd4809; ROM2[7235]<=16'd0; ROM3[7235]<=16'd23769; ROM4[7235]<=16'd57268;
ROM1[7236]<=16'd4795; ROM2[7236]<=16'd0; ROM3[7236]<=16'd23773; ROM4[7236]<=16'd57268;
ROM1[7237]<=16'd4774; ROM2[7237]<=16'd0; ROM3[7237]<=16'd23765; ROM4[7237]<=16'd57257;
ROM1[7238]<=16'd4769; ROM2[7238]<=16'd0; ROM3[7238]<=16'd23752; ROM4[7238]<=16'd57246;
ROM1[7239]<=16'd4820; ROM2[7239]<=16'd0; ROM3[7239]<=16'd23757; ROM4[7239]<=16'd57265;
ROM1[7240]<=16'd4868; ROM2[7240]<=16'd0; ROM3[7240]<=16'd23771; ROM4[7240]<=16'd57290;
ROM1[7241]<=16'd4842; ROM2[7241]<=16'd0; ROM3[7241]<=16'd23758; ROM4[7241]<=16'd57274;
ROM1[7242]<=16'd4825; ROM2[7242]<=16'd0; ROM3[7242]<=16'd23765; ROM4[7242]<=16'd57277;
ROM1[7243]<=16'd4804; ROM2[7243]<=16'd0; ROM3[7243]<=16'd23770; ROM4[7243]<=16'd57278;
ROM1[7244]<=16'd4781; ROM2[7244]<=16'd0; ROM3[7244]<=16'd23767; ROM4[7244]<=16'd57267;
ROM1[7245]<=16'd4782; ROM2[7245]<=16'd0; ROM3[7245]<=16'd23788; ROM4[7245]<=16'd57282;
ROM1[7246]<=16'd4790; ROM2[7246]<=16'd0; ROM3[7246]<=16'd23803; ROM4[7246]<=16'd57296;
ROM1[7247]<=16'd4795; ROM2[7247]<=16'd0; ROM3[7247]<=16'd23783; ROM4[7247]<=16'd57282;
ROM1[7248]<=16'd4810; ROM2[7248]<=16'd0; ROM3[7248]<=16'd23754; ROM4[7248]<=16'd57266;
ROM1[7249]<=16'd4839; ROM2[7249]<=16'd0; ROM3[7249]<=16'd23766; ROM4[7249]<=16'd57283;
ROM1[7250]<=16'd4840; ROM2[7250]<=16'd0; ROM3[7250]<=16'd23781; ROM4[7250]<=16'd57294;
ROM1[7251]<=16'd4814; ROM2[7251]<=16'd0; ROM3[7251]<=16'd23786; ROM4[7251]<=16'd57289;
ROM1[7252]<=16'd4788; ROM2[7252]<=16'd0; ROM3[7252]<=16'd23782; ROM4[7252]<=16'd57281;
ROM1[7253]<=16'd4772; ROM2[7253]<=16'd0; ROM3[7253]<=16'd23780; ROM4[7253]<=16'd57273;
ROM1[7254]<=16'd4765; ROM2[7254]<=16'd0; ROM3[7254]<=16'd23773; ROM4[7254]<=16'd57265;
ROM1[7255]<=16'd4783; ROM2[7255]<=16'd0; ROM3[7255]<=16'd23773; ROM4[7255]<=16'd57266;
ROM1[7256]<=16'd4826; ROM2[7256]<=16'd0; ROM3[7256]<=16'd23772; ROM4[7256]<=16'd57274;
ROM1[7257]<=16'd4841; ROM2[7257]<=16'd0; ROM3[7257]<=16'd23759; ROM4[7257]<=16'd57273;
ROM1[7258]<=16'd4823; ROM2[7258]<=16'd0; ROM3[7258]<=16'd23753; ROM4[7258]<=16'd57265;
ROM1[7259]<=16'd4802; ROM2[7259]<=16'd0; ROM3[7259]<=16'd23762; ROM4[7259]<=16'd57261;
ROM1[7260]<=16'd4799; ROM2[7260]<=16'd0; ROM3[7260]<=16'd23785; ROM4[7260]<=16'd57269;
ROM1[7261]<=16'd4788; ROM2[7261]<=16'd0; ROM3[7261]<=16'd23793; ROM4[7261]<=16'd57274;
ROM1[7262]<=16'd4774; ROM2[7262]<=16'd0; ROM3[7262]<=16'd23791; ROM4[7262]<=16'd57266;
ROM1[7263]<=16'd4788; ROM2[7263]<=16'd0; ROM3[7263]<=16'd23793; ROM4[7263]<=16'd57273;
ROM1[7264]<=16'd4818; ROM2[7264]<=16'd0; ROM3[7264]<=16'd23789; ROM4[7264]<=16'd57279;
ROM1[7265]<=16'd4852; ROM2[7265]<=16'd0; ROM3[7265]<=16'd23788; ROM4[7265]<=16'd57284;
ROM1[7266]<=16'd4852; ROM2[7266]<=16'd0; ROM3[7266]<=16'd23792; ROM4[7266]<=16'd57292;
ROM1[7267]<=16'd4830; ROM2[7267]<=16'd0; ROM3[7267]<=16'd23791; ROM4[7267]<=16'd57290;
ROM1[7268]<=16'd4820; ROM2[7268]<=16'd0; ROM3[7268]<=16'd23805; ROM4[7268]<=16'd57300;
ROM1[7269]<=16'd4825; ROM2[7269]<=16'd0; ROM3[7269]<=16'd23820; ROM4[7269]<=16'd57315;
ROM1[7270]<=16'd4818; ROM2[7270]<=16'd0; ROM3[7270]<=16'd23819; ROM4[7270]<=16'd57315;
ROM1[7271]<=16'd4827; ROM2[7271]<=16'd0; ROM3[7271]<=16'd23822; ROM4[7271]<=16'd57323;
ROM1[7272]<=16'd4842; ROM2[7272]<=16'd0; ROM3[7272]<=16'd23807; ROM4[7272]<=16'd57316;
ROM1[7273]<=16'd4849; ROM2[7273]<=16'd0; ROM3[7273]<=16'd23771; ROM4[7273]<=16'd57293;
ROM1[7274]<=16'd4849; ROM2[7274]<=16'd0; ROM3[7274]<=16'd23761; ROM4[7274]<=16'd57282;
ROM1[7275]<=16'd4842; ROM2[7275]<=16'd0; ROM3[7275]<=16'd23773; ROM4[7275]<=16'd57286;
ROM1[7276]<=16'd4826; ROM2[7276]<=16'd0; ROM3[7276]<=16'd23788; ROM4[7276]<=16'd57291;
ROM1[7277]<=16'd4797; ROM2[7277]<=16'd0; ROM3[7277]<=16'd23782; ROM4[7277]<=16'd57279;
ROM1[7278]<=16'd4788; ROM2[7278]<=16'd0; ROM3[7278]<=16'd23785; ROM4[7278]<=16'd57278;
ROM1[7279]<=16'd4778; ROM2[7279]<=16'd0; ROM3[7279]<=16'd23778; ROM4[7279]<=16'd57271;
ROM1[7280]<=16'd4777; ROM2[7280]<=16'd0; ROM3[7280]<=16'd23754; ROM4[7280]<=16'd57254;
ROM1[7281]<=16'd4818; ROM2[7281]<=16'd0; ROM3[7281]<=16'd23756; ROM4[7281]<=16'd57263;
ROM1[7282]<=16'd4854; ROM2[7282]<=16'd0; ROM3[7282]<=16'd23772; ROM4[7282]<=16'd57283;
ROM1[7283]<=16'd4850; ROM2[7283]<=16'd0; ROM3[7283]<=16'd23775; ROM4[7283]<=16'd57283;
ROM1[7284]<=16'd4825; ROM2[7284]<=16'd0; ROM3[7284]<=16'd23772; ROM4[7284]<=16'd57273;
ROM1[7285]<=16'd4810; ROM2[7285]<=16'd0; ROM3[7285]<=16'd23782; ROM4[7285]<=16'd57277;
ROM1[7286]<=16'd4792; ROM2[7286]<=16'd0; ROM3[7286]<=16'd23782; ROM4[7286]<=16'd57274;
ROM1[7287]<=16'd4782; ROM2[7287]<=16'd0; ROM3[7287]<=16'd23782; ROM4[7287]<=16'd57272;
ROM1[7288]<=16'd4801; ROM2[7288]<=16'd0; ROM3[7288]<=16'd23790; ROM4[7288]<=16'd57281;
ROM1[7289]<=16'd4832; ROM2[7289]<=16'd0; ROM3[7289]<=16'd23788; ROM4[7289]<=16'd57286;
ROM1[7290]<=16'd4848; ROM2[7290]<=16'd0; ROM3[7290]<=16'd23771; ROM4[7290]<=16'd57276;
ROM1[7291]<=16'd4836; ROM2[7291]<=16'd0; ROM3[7291]<=16'd23766; ROM4[7291]<=16'd57272;
ROM1[7292]<=16'd4833; ROM2[7292]<=16'd0; ROM3[7292]<=16'd23786; ROM4[7292]<=16'd57287;
ROM1[7293]<=16'd4823; ROM2[7293]<=16'd0; ROM3[7293]<=16'd23798; ROM4[7293]<=16'd57293;
ROM1[7294]<=16'd4810; ROM2[7294]<=16'd0; ROM3[7294]<=16'd23799; ROM4[7294]<=16'd57293;
ROM1[7295]<=16'd4797; ROM2[7295]<=16'd0; ROM3[7295]<=16'd23803; ROM4[7295]<=16'd57293;
ROM1[7296]<=16'd4791; ROM2[7296]<=16'd0; ROM3[7296]<=16'd23798; ROM4[7296]<=16'd57286;
ROM1[7297]<=16'd4807; ROM2[7297]<=16'd0; ROM3[7297]<=16'd23785; ROM4[7297]<=16'd57282;
ROM1[7298]<=16'd4847; ROM2[7298]<=16'd0; ROM3[7298]<=16'd23784; ROM4[7298]<=16'd57293;
ROM1[7299]<=16'd4864; ROM2[7299]<=16'd0; ROM3[7299]<=16'd23794; ROM4[7299]<=16'd57300;
ROM1[7300]<=16'd4847; ROM2[7300]<=16'd0; ROM3[7300]<=16'd23793; ROM4[7300]<=16'd57299;
ROM1[7301]<=16'd4821; ROM2[7301]<=16'd0; ROM3[7301]<=16'd23791; ROM4[7301]<=16'd57291;
ROM1[7302]<=16'd4795; ROM2[7302]<=16'd0; ROM3[7302]<=16'd23789; ROM4[7302]<=16'd57279;
ROM1[7303]<=16'd4770; ROM2[7303]<=16'd0; ROM3[7303]<=16'd23783; ROM4[7303]<=16'd57268;
ROM1[7304]<=16'd4771; ROM2[7304]<=16'd0; ROM3[7304]<=16'd23791; ROM4[7304]<=16'd57273;
ROM1[7305]<=16'd4800; ROM2[7305]<=16'd0; ROM3[7305]<=16'd23800; ROM4[7305]<=16'd57286;
ROM1[7306]<=16'd4826; ROM2[7306]<=16'd0; ROM3[7306]<=16'd23786; ROM4[7306]<=16'd57281;
ROM1[7307]<=16'd4843; ROM2[7307]<=16'd0; ROM3[7307]<=16'd23778; ROM4[7307]<=16'd57279;
ROM1[7308]<=16'd4852; ROM2[7308]<=16'd0; ROM3[7308]<=16'd23798; ROM4[7308]<=16'd57297;
ROM1[7309]<=16'd4829; ROM2[7309]<=16'd0; ROM3[7309]<=16'd23801; ROM4[7309]<=16'd57295;
ROM1[7310]<=16'd4797; ROM2[7310]<=16'd0; ROM3[7310]<=16'd23792; ROM4[7310]<=16'd57279;
ROM1[7311]<=16'd4785; ROM2[7311]<=16'd0; ROM3[7311]<=16'd23800; ROM4[7311]<=16'd57284;
ROM1[7312]<=16'd4772; ROM2[7312]<=16'd0; ROM3[7312]<=16'd23797; ROM4[7312]<=16'd57280;
ROM1[7313]<=16'd4786; ROM2[7313]<=16'd0; ROM3[7313]<=16'd23799; ROM4[7313]<=16'd57281;
ROM1[7314]<=16'd4829; ROM2[7314]<=16'd0; ROM3[7314]<=16'd23807; ROM4[7314]<=16'd57297;
ROM1[7315]<=16'd4853; ROM2[7315]<=16'd0; ROM3[7315]<=16'd23789; ROM4[7315]<=16'd57294;
ROM1[7316]<=16'd4851; ROM2[7316]<=16'd0; ROM3[7316]<=16'd23787; ROM4[7316]<=16'd57291;
ROM1[7317]<=16'd4839; ROM2[7317]<=16'd0; ROM3[7317]<=16'd23795; ROM4[7317]<=16'd57293;
ROM1[7318]<=16'd4814; ROM2[7318]<=16'd0; ROM3[7318]<=16'd23787; ROM4[7318]<=16'd57283;
ROM1[7319]<=16'd4806; ROM2[7319]<=16'd0; ROM3[7319]<=16'd23797; ROM4[7319]<=16'd57286;
ROM1[7320]<=16'd4785; ROM2[7320]<=16'd0; ROM3[7320]<=16'd23799; ROM4[7320]<=16'd57281;
ROM1[7321]<=16'd4771; ROM2[7321]<=16'd0; ROM3[7321]<=16'd23783; ROM4[7321]<=16'd57272;
ROM1[7322]<=16'd4803; ROM2[7322]<=16'd0; ROM3[7322]<=16'd23786; ROM4[7322]<=16'd57280;
ROM1[7323]<=16'd4837; ROM2[7323]<=16'd0; ROM3[7323]<=16'd23777; ROM4[7323]<=16'd57282;
ROM1[7324]<=16'd4842; ROM2[7324]<=16'd0; ROM3[7324]<=16'd23766; ROM4[7324]<=16'd57278;
ROM1[7325]<=16'd4842; ROM2[7325]<=16'd0; ROM3[7325]<=16'd23783; ROM4[7325]<=16'd57291;
ROM1[7326]<=16'd4831; ROM2[7326]<=16'd0; ROM3[7326]<=16'd23805; ROM4[7326]<=16'd57305;
ROM1[7327]<=16'd4804; ROM2[7327]<=16'd0; ROM3[7327]<=16'd23795; ROM4[7327]<=16'd57293;
ROM1[7328]<=16'd4782; ROM2[7328]<=16'd0; ROM3[7328]<=16'd23787; ROM4[7328]<=16'd57282;
ROM1[7329]<=16'd4766; ROM2[7329]<=16'd0; ROM3[7329]<=16'd23779; ROM4[7329]<=16'd57269;
ROM1[7330]<=16'd4773; ROM2[7330]<=16'd0; ROM3[7330]<=16'd23769; ROM4[7330]<=16'd57266;
ROM1[7331]<=16'd4809; ROM2[7331]<=16'd0; ROM3[7331]<=16'd23767; ROM4[7331]<=16'd57276;
ROM1[7332]<=16'd4838; ROM2[7332]<=16'd0; ROM3[7332]<=16'd23777; ROM4[7332]<=16'd57288;
ROM1[7333]<=16'd4835; ROM2[7333]<=16'd0; ROM3[7333]<=16'd23780; ROM4[7333]<=16'd57292;
ROM1[7334]<=16'd4800; ROM2[7334]<=16'd0; ROM3[7334]<=16'd23764; ROM4[7334]<=16'd57272;
ROM1[7335]<=16'd4778; ROM2[7335]<=16'd0; ROM3[7335]<=16'd23761; ROM4[7335]<=16'd57262;
ROM1[7336]<=16'd4773; ROM2[7336]<=16'd0; ROM3[7336]<=16'd23765; ROM4[7336]<=16'd57263;
ROM1[7337]<=16'd4776; ROM2[7337]<=16'd0; ROM3[7337]<=16'd23779; ROM4[7337]<=16'd57272;
ROM1[7338]<=16'd4794; ROM2[7338]<=16'd0; ROM3[7338]<=16'd23785; ROM4[7338]<=16'd57281;
ROM1[7339]<=16'd4815; ROM2[7339]<=16'd0; ROM3[7339]<=16'd23764; ROM4[7339]<=16'd57273;
ROM1[7340]<=16'd4829; ROM2[7340]<=16'd0; ROM3[7340]<=16'd23747; ROM4[7340]<=16'd57265;
ROM1[7341]<=16'd4821; ROM2[7341]<=16'd0; ROM3[7341]<=16'd23742; ROM4[7341]<=16'd57259;
ROM1[7342]<=16'd4813; ROM2[7342]<=16'd0; ROM3[7342]<=16'd23751; ROM4[7342]<=16'd57263;
ROM1[7343]<=16'd4798; ROM2[7343]<=16'd0; ROM3[7343]<=16'd23764; ROM4[7343]<=16'd57267;
ROM1[7344]<=16'd4778; ROM2[7344]<=16'd0; ROM3[7344]<=16'd23767; ROM4[7344]<=16'd57267;
ROM1[7345]<=16'd4776; ROM2[7345]<=16'd0; ROM3[7345]<=16'd23778; ROM4[7345]<=16'd57276;
ROM1[7346]<=16'd4781; ROM2[7346]<=16'd0; ROM3[7346]<=16'd23781; ROM4[7346]<=16'd57276;
ROM1[7347]<=16'd4799; ROM2[7347]<=16'd0; ROM3[7347]<=16'd23772; ROM4[7347]<=16'd57271;
ROM1[7348]<=16'd4815; ROM2[7348]<=16'd0; ROM3[7348]<=16'd23744; ROM4[7348]<=16'd57253;
ROM1[7349]<=16'd4810; ROM2[7349]<=16'd0; ROM3[7349]<=16'd23731; ROM4[7349]<=16'd57243;
ROM1[7350]<=16'd4801; ROM2[7350]<=16'd0; ROM3[7350]<=16'd23744; ROM4[7350]<=16'd57252;
ROM1[7351]<=16'd4791; ROM2[7351]<=16'd0; ROM3[7351]<=16'd23758; ROM4[7351]<=16'd57261;
ROM1[7352]<=16'd4786; ROM2[7352]<=16'd0; ROM3[7352]<=16'd23774; ROM4[7352]<=16'd57271;
ROM1[7353]<=16'd4772; ROM2[7353]<=16'd0; ROM3[7353]<=16'd23783; ROM4[7353]<=16'd57271;
ROM1[7354]<=16'd4772; ROM2[7354]<=16'd0; ROM3[7354]<=16'd23792; ROM4[7354]<=16'd57281;
ROM1[7355]<=16'd4785; ROM2[7355]<=16'd0; ROM3[7355]<=16'd23787; ROM4[7355]<=16'd57284;
ROM1[7356]<=16'd4819; ROM2[7356]<=16'd0; ROM3[7356]<=16'd23770; ROM4[7356]<=16'd57281;
ROM1[7357]<=16'd4841; ROM2[7357]<=16'd0; ROM3[7357]<=16'd23766; ROM4[7357]<=16'd57287;
ROM1[7358]<=16'd4835; ROM2[7358]<=16'd0; ROM3[7358]<=16'd23776; ROM4[7358]<=16'd57290;
ROM1[7359]<=16'd4823; ROM2[7359]<=16'd0; ROM3[7359]<=16'd23784; ROM4[7359]<=16'd57288;
ROM1[7360]<=16'd4808; ROM2[7360]<=16'd0; ROM3[7360]<=16'd23790; ROM4[7360]<=16'd57291;
ROM1[7361]<=16'd4789; ROM2[7361]<=16'd0; ROM3[7361]<=16'd23790; ROM4[7361]<=16'd57286;
ROM1[7362]<=16'd4769; ROM2[7362]<=16'd0; ROM3[7362]<=16'd23778; ROM4[7362]<=16'd57275;
ROM1[7363]<=16'd4780; ROM2[7363]<=16'd0; ROM3[7363]<=16'd23776; ROM4[7363]<=16'd57279;
ROM1[7364]<=16'd4817; ROM2[7364]<=16'd0; ROM3[7364]<=16'd23778; ROM4[7364]<=16'd57285;
ROM1[7365]<=16'd4842; ROM2[7365]<=16'd0; ROM3[7365]<=16'd23766; ROM4[7365]<=16'd57281;
ROM1[7366]<=16'd4837; ROM2[7366]<=16'd0; ROM3[7366]<=16'd23759; ROM4[7366]<=16'd57276;
ROM1[7367]<=16'd4825; ROM2[7367]<=16'd0; ROM3[7367]<=16'd23770; ROM4[7367]<=16'd57284;
ROM1[7368]<=16'd4811; ROM2[7368]<=16'd0; ROM3[7368]<=16'd23782; ROM4[7368]<=16'd57289;
ROM1[7369]<=16'd4808; ROM2[7369]<=16'd0; ROM3[7369]<=16'd23793; ROM4[7369]<=16'd57295;
ROM1[7370]<=16'd4802; ROM2[7370]<=16'd0; ROM3[7370]<=16'd23798; ROM4[7370]<=16'd57296;
ROM1[7371]<=16'd4800; ROM2[7371]<=16'd0; ROM3[7371]<=16'd23795; ROM4[7371]<=16'd57289;
ROM1[7372]<=16'd4824; ROM2[7372]<=16'd0; ROM3[7372]<=16'd23790; ROM4[7372]<=16'd57289;
ROM1[7373]<=16'd4857; ROM2[7373]<=16'd0; ROM3[7373]<=16'd23774; ROM4[7373]<=16'd57289;
ROM1[7374]<=16'd4865; ROM2[7374]<=16'd0; ROM3[7374]<=16'd23774; ROM4[7374]<=16'd57291;
ROM1[7375]<=16'd4849; ROM2[7375]<=16'd0; ROM3[7375]<=16'd23779; ROM4[7375]<=16'd57295;
ROM1[7376]<=16'd4815; ROM2[7376]<=16'd0; ROM3[7376]<=16'd23774; ROM4[7376]<=16'd57287;
ROM1[7377]<=16'd4794; ROM2[7377]<=16'd0; ROM3[7377]<=16'd23779; ROM4[7377]<=16'd57280;
ROM1[7378]<=16'd4782; ROM2[7378]<=16'd0; ROM3[7378]<=16'd23789; ROM4[7378]<=16'd57285;
ROM1[7379]<=16'd4777; ROM2[7379]<=16'd0; ROM3[7379]<=16'd23784; ROM4[7379]<=16'd57279;
ROM1[7380]<=16'd4778; ROM2[7380]<=16'd0; ROM3[7380]<=16'd23759; ROM4[7380]<=16'd57264;
ROM1[7381]<=16'd4802; ROM2[7381]<=16'd0; ROM3[7381]<=16'd23743; ROM4[7381]<=16'd57262;
ROM1[7382]<=16'd4824; ROM2[7382]<=16'd0; ROM3[7382]<=16'd23737; ROM4[7382]<=16'd57262;
ROM1[7383]<=16'd4818; ROM2[7383]<=16'd0; ROM3[7383]<=16'd23743; ROM4[7383]<=16'd57265;
ROM1[7384]<=16'd4798; ROM2[7384]<=16'd0; ROM3[7384]<=16'd23750; ROM4[7384]<=16'd57262;
ROM1[7385]<=16'd4773; ROM2[7385]<=16'd0; ROM3[7385]<=16'd23750; ROM4[7385]<=16'd57256;
ROM1[7386]<=16'd4770; ROM2[7386]<=16'd0; ROM3[7386]<=16'd23763; ROM4[7386]<=16'd57266;
ROM1[7387]<=16'd4773; ROM2[7387]<=16'd0; ROM3[7387]<=16'd23780; ROM4[7387]<=16'd57275;
ROM1[7388]<=16'd4783; ROM2[7388]<=16'd0; ROM3[7388]<=16'd23779; ROM4[7388]<=16'd57277;
ROM1[7389]<=16'd4789; ROM2[7389]<=16'd0; ROM3[7389]<=16'd23743; ROM4[7389]<=16'd57255;
ROM1[7390]<=16'd4801; ROM2[7390]<=16'd0; ROM3[7390]<=16'd23715; ROM4[7390]<=16'd57237;
ROM1[7391]<=16'd4800; ROM2[7391]<=16'd0; ROM3[7391]<=16'd23714; ROM4[7391]<=16'd57237;
ROM1[7392]<=16'd4796; ROM2[7392]<=16'd0; ROM3[7392]<=16'd23731; ROM4[7392]<=16'd57250;
ROM1[7393]<=16'd4803; ROM2[7393]<=16'd0; ROM3[7393]<=16'd23761; ROM4[7393]<=16'd57270;
ROM1[7394]<=16'd4786; ROM2[7394]<=16'd0; ROM3[7394]<=16'd23766; ROM4[7394]<=16'd57273;
ROM1[7395]<=16'd4769; ROM2[7395]<=16'd0; ROM3[7395]<=16'd23769; ROM4[7395]<=16'd57272;
ROM1[7396]<=16'd4790; ROM2[7396]<=16'd0; ROM3[7396]<=16'd23778; ROM4[7396]<=16'd57285;
ROM1[7397]<=16'd4817; ROM2[7397]<=16'd0; ROM3[7397]<=16'd23768; ROM4[7397]<=16'd57286;
ROM1[7398]<=16'd4832; ROM2[7398]<=16'd0; ROM3[7398]<=16'd23747; ROM4[7398]<=16'd57275;
ROM1[7399]<=16'd4839; ROM2[7399]<=16'd0; ROM3[7399]<=16'd23740; ROM4[7399]<=16'd57273;
ROM1[7400]<=16'd4826; ROM2[7400]<=16'd0; ROM3[7400]<=16'd23742; ROM4[7400]<=16'd57272;
ROM1[7401]<=16'd4814; ROM2[7401]<=16'd0; ROM3[7401]<=16'd23757; ROM4[7401]<=16'd57279;
ROM1[7402]<=16'd4814; ROM2[7402]<=16'd0; ROM3[7402]<=16'd23777; ROM4[7402]<=16'd57292;
ROM1[7403]<=16'd4795; ROM2[7403]<=16'd0; ROM3[7403]<=16'd23781; ROM4[7403]<=16'd57290;
ROM1[7404]<=16'd4790; ROM2[7404]<=16'd0; ROM3[7404]<=16'd23783; ROM4[7404]<=16'd57290;
ROM1[7405]<=16'd4806; ROM2[7405]<=16'd0; ROM3[7405]<=16'd23783; ROM4[7405]<=16'd57292;
ROM1[7406]<=16'd4829; ROM2[7406]<=16'd0; ROM3[7406]<=16'd23760; ROM4[7406]<=16'd57275;
ROM1[7407]<=16'd4835; ROM2[7407]<=16'd0; ROM3[7407]<=16'd23745; ROM4[7407]<=16'd57266;
ROM1[7408]<=16'd4832; ROM2[7408]<=16'd0; ROM3[7408]<=16'd23757; ROM4[7408]<=16'd57278;
ROM1[7409]<=16'd4822; ROM2[7409]<=16'd0; ROM3[7409]<=16'd23774; ROM4[7409]<=16'd57286;
ROM1[7410]<=16'd4809; ROM2[7410]<=16'd0; ROM3[7410]<=16'd23787; ROM4[7410]<=16'd57294;
ROM1[7411]<=16'd4809; ROM2[7411]<=16'd0; ROM3[7411]<=16'd23814; ROM4[7411]<=16'd57309;
ROM1[7412]<=16'd4815; ROM2[7412]<=16'd0; ROM3[7412]<=16'd23837; ROM4[7412]<=16'd57328;
ROM1[7413]<=16'd4815; ROM2[7413]<=16'd0; ROM3[7413]<=16'd23828; ROM4[7413]<=16'd57326;
ROM1[7414]<=16'd4834; ROM2[7414]<=16'd0; ROM3[7414]<=16'd23808; ROM4[7414]<=16'd57314;
ROM1[7415]<=16'd4863; ROM2[7415]<=16'd0; ROM3[7415]<=16'd23791; ROM4[7415]<=16'd57310;
ROM1[7416]<=16'd4855; ROM2[7416]<=16'd0; ROM3[7416]<=16'd23782; ROM4[7416]<=16'd57301;
ROM1[7417]<=16'd4845; ROM2[7417]<=16'd0; ROM3[7417]<=16'd23801; ROM4[7417]<=16'd57308;
ROM1[7418]<=16'd4834; ROM2[7418]<=16'd0; ROM3[7418]<=16'd23813; ROM4[7418]<=16'd57315;
ROM1[7419]<=16'd4805; ROM2[7419]<=16'd0; ROM3[7419]<=16'd23800; ROM4[7419]<=16'd57301;
ROM1[7420]<=16'd4784; ROM2[7420]<=16'd0; ROM3[7420]<=16'd23792; ROM4[7420]<=16'd57286;
ROM1[7421]<=16'd4785; ROM2[7421]<=16'd0; ROM3[7421]<=16'd23783; ROM4[7421]<=16'd57278;
ROM1[7422]<=16'd4808; ROM2[7422]<=16'd0; ROM3[7422]<=16'd23776; ROM4[7422]<=16'd57278;
ROM1[7423]<=16'd4844; ROM2[7423]<=16'd0; ROM3[7423]<=16'd23767; ROM4[7423]<=16'd57282;
ROM1[7424]<=16'd4848; ROM2[7424]<=16'd0; ROM3[7424]<=16'd23760; ROM4[7424]<=16'd57281;
ROM1[7425]<=16'd4830; ROM2[7425]<=16'd0; ROM3[7425]<=16'd23756; ROM4[7425]<=16'd57276;
ROM1[7426]<=16'd4811; ROM2[7426]<=16'd0; ROM3[7426]<=16'd23760; ROM4[7426]<=16'd57276;
ROM1[7427]<=16'd4804; ROM2[7427]<=16'd0; ROM3[7427]<=16'd23769; ROM4[7427]<=16'd57279;
ROM1[7428]<=16'd4790; ROM2[7428]<=16'd0; ROM3[7428]<=16'd23768; ROM4[7428]<=16'd57271;
ROM1[7429]<=16'd4787; ROM2[7429]<=16'd0; ROM3[7429]<=16'd23767; ROM4[7429]<=16'd57271;
ROM1[7430]<=16'd4806; ROM2[7430]<=16'd0; ROM3[7430]<=16'd23762; ROM4[7430]<=16'd57271;
ROM1[7431]<=16'd4832; ROM2[7431]<=16'd0; ROM3[7431]<=16'd23738; ROM4[7431]<=16'd57261;
ROM1[7432]<=16'd4855; ROM2[7432]<=16'd0; ROM3[7432]<=16'd23737; ROM4[7432]<=16'd57269;
ROM1[7433]<=16'd4852; ROM2[7433]<=16'd0; ROM3[7433]<=16'd23746; ROM4[7433]<=16'd57276;
ROM1[7434]<=16'd4833; ROM2[7434]<=16'd0; ROM3[7434]<=16'd23748; ROM4[7434]<=16'd57276;
ROM1[7435]<=16'd4805; ROM2[7435]<=16'd0; ROM3[7435]<=16'd23742; ROM4[7435]<=16'd57263;
ROM1[7436]<=16'd4767; ROM2[7436]<=16'd0; ROM3[7436]<=16'd23730; ROM4[7436]<=16'd57245;
ROM1[7437]<=16'd4754; ROM2[7437]<=16'd0; ROM3[7437]<=16'd23729; ROM4[7437]<=16'd57239;
ROM1[7438]<=16'd4772; ROM2[7438]<=16'd0; ROM3[7438]<=16'd23729; ROM4[7438]<=16'd57240;
ROM1[7439]<=16'd4805; ROM2[7439]<=16'd0; ROM3[7439]<=16'd23723; ROM4[7439]<=16'd57245;
ROM1[7440]<=16'd4836; ROM2[7440]<=16'd0; ROM3[7440]<=16'd23717; ROM4[7440]<=16'd57245;
ROM1[7441]<=16'd4844; ROM2[7441]<=16'd0; ROM3[7441]<=16'd23727; ROM4[7441]<=16'd57255;
ROM1[7442]<=16'd4834; ROM2[7442]<=16'd0; ROM3[7442]<=16'd23743; ROM4[7442]<=16'd57263;
ROM1[7443]<=16'd4828; ROM2[7443]<=16'd0; ROM3[7443]<=16'd23771; ROM4[7443]<=16'd57275;
ROM1[7444]<=16'd4815; ROM2[7444]<=16'd0; ROM3[7444]<=16'd23777; ROM4[7444]<=16'd57281;
ROM1[7445]<=16'd4774; ROM2[7445]<=16'd0; ROM3[7445]<=16'd23754; ROM4[7445]<=16'd57255;
ROM1[7446]<=16'd4763; ROM2[7446]<=16'd0; ROM3[7446]<=16'd23745; ROM4[7446]<=16'd57244;
ROM1[7447]<=16'd4787; ROM2[7447]<=16'd0; ROM3[7447]<=16'd23744; ROM4[7447]<=16'd57252;
ROM1[7448]<=16'd4819; ROM2[7448]<=16'd0; ROM3[7448]<=16'd23733; ROM4[7448]<=16'd57255;
ROM1[7449]<=16'd4838; ROM2[7449]<=16'd0; ROM3[7449]<=16'd23743; ROM4[7449]<=16'd57267;
ROM1[7450]<=16'd4844; ROM2[7450]<=16'd0; ROM3[7450]<=16'd23770; ROM4[7450]<=16'd57289;
ROM1[7451]<=16'd4827; ROM2[7451]<=16'd0; ROM3[7451]<=16'd23778; ROM4[7451]<=16'd57290;
ROM1[7452]<=16'd4812; ROM2[7452]<=16'd0; ROM3[7452]<=16'd23783; ROM4[7452]<=16'd57288;
ROM1[7453]<=16'd4802; ROM2[7453]<=16'd0; ROM3[7453]<=16'd23793; ROM4[7453]<=16'd57292;
ROM1[7454]<=16'd4790; ROM2[7454]<=16'd0; ROM3[7454]<=16'd23784; ROM4[7454]<=16'd57285;
ROM1[7455]<=16'd4803; ROM2[7455]<=16'd0; ROM3[7455]<=16'd23776; ROM4[7455]<=16'd57287;
ROM1[7456]<=16'd4835; ROM2[7456]<=16'd0; ROM3[7456]<=16'd23769; ROM4[7456]<=16'd57287;
ROM1[7457]<=16'd4849; ROM2[7457]<=16'd0; ROM3[7457]<=16'd23761; ROM4[7457]<=16'd57288;
ROM1[7458]<=16'd4841; ROM2[7458]<=16'd0; ROM3[7458]<=16'd23767; ROM4[7458]<=16'd57290;
ROM1[7459]<=16'd4821; ROM2[7459]<=16'd0; ROM3[7459]<=16'd23774; ROM4[7459]<=16'd57285;
ROM1[7460]<=16'd4807; ROM2[7460]<=16'd0; ROM3[7460]<=16'd23782; ROM4[7460]<=16'd57288;
ROM1[7461]<=16'd4794; ROM2[7461]<=16'd0; ROM3[7461]<=16'd23786; ROM4[7461]<=16'd57286;
ROM1[7462]<=16'd4780; ROM2[7462]<=16'd0; ROM3[7462]<=16'd23786; ROM4[7462]<=16'd57282;
ROM1[7463]<=16'd4787; ROM2[7463]<=16'd0; ROM3[7463]<=16'd23785; ROM4[7463]<=16'd57279;
ROM1[7464]<=16'd4823; ROM2[7464]<=16'd0; ROM3[7464]<=16'd23780; ROM4[7464]<=16'd57280;
ROM1[7465]<=16'd4851; ROM2[7465]<=16'd0; ROM3[7465]<=16'd23770; ROM4[7465]<=16'd57283;
ROM1[7466]<=16'd4844; ROM2[7466]<=16'd0; ROM3[7466]<=16'd23766; ROM4[7466]<=16'd57276;
ROM1[7467]<=16'd4827; ROM2[7467]<=16'd0; ROM3[7467]<=16'd23771; ROM4[7467]<=16'd57275;
ROM1[7468]<=16'd4804; ROM2[7468]<=16'd0; ROM3[7468]<=16'd23777; ROM4[7468]<=16'd57272;
ROM1[7469]<=16'd4807; ROM2[7469]<=16'd0; ROM3[7469]<=16'd23797; ROM4[7469]<=16'd57287;
ROM1[7470]<=16'd4816; ROM2[7470]<=16'd0; ROM3[7470]<=16'd23821; ROM4[7470]<=16'd57310;
ROM1[7471]<=16'd4796; ROM2[7471]<=16'd0; ROM3[7471]<=16'd23799; ROM4[7471]<=16'd57287;
ROM1[7472]<=16'd4803; ROM2[7472]<=16'd0; ROM3[7472]<=16'd23774; ROM4[7472]<=16'd57268;
ROM1[7473]<=16'd4822; ROM2[7473]<=16'd0; ROM3[7473]<=16'd23753; ROM4[7473]<=16'd57260;
ROM1[7474]<=16'd4816; ROM2[7474]<=16'd0; ROM3[7474]<=16'd23744; ROM4[7474]<=16'd57256;
ROM1[7475]<=16'd4823; ROM2[7475]<=16'd0; ROM3[7475]<=16'd23763; ROM4[7475]<=16'd57271;
ROM1[7476]<=16'd4811; ROM2[7476]<=16'd0; ROM3[7476]<=16'd23776; ROM4[7476]<=16'd57280;
ROM1[7477]<=16'd4788; ROM2[7477]<=16'd0; ROM3[7477]<=16'd23772; ROM4[7477]<=16'd57275;
ROM1[7478]<=16'd4769; ROM2[7478]<=16'd0; ROM3[7478]<=16'd23766; ROM4[7478]<=16'd57266;
ROM1[7479]<=16'd4766; ROM2[7479]<=16'd0; ROM3[7479]<=16'd23763; ROM4[7479]<=16'd57265;
ROM1[7480]<=16'd4784; ROM2[7480]<=16'd0; ROM3[7480]<=16'd23760; ROM4[7480]<=16'd57262;
ROM1[7481]<=16'd4815; ROM2[7481]<=16'd0; ROM3[7481]<=16'd23745; ROM4[7481]<=16'd57256;
ROM1[7482]<=16'd4827; ROM2[7482]<=16'd0; ROM3[7482]<=16'd23732; ROM4[7482]<=16'd57251;
ROM1[7483]<=16'd4820; ROM2[7483]<=16'd0; ROM3[7483]<=16'd23737; ROM4[7483]<=16'd57259;
ROM1[7484]<=16'd4808; ROM2[7484]<=16'd0; ROM3[7484]<=16'd23752; ROM4[7484]<=16'd57269;
ROM1[7485]<=16'd4802; ROM2[7485]<=16'd0; ROM3[7485]<=16'd23768; ROM4[7485]<=16'd57279;
ROM1[7486]<=16'd4789; ROM2[7486]<=16'd0; ROM3[7486]<=16'd23770; ROM4[7486]<=16'd57278;
ROM1[7487]<=16'd4791; ROM2[7487]<=16'd0; ROM3[7487]<=16'd23779; ROM4[7487]<=16'd57280;
ROM1[7488]<=16'd4808; ROM2[7488]<=16'd0; ROM3[7488]<=16'd23782; ROM4[7488]<=16'd57283;
ROM1[7489]<=16'd4816; ROM2[7489]<=16'd0; ROM3[7489]<=16'd23752; ROM4[7489]<=16'd57260;
ROM1[7490]<=16'd4828; ROM2[7490]<=16'd0; ROM3[7490]<=16'd23734; ROM4[7490]<=16'd57248;
ROM1[7491]<=16'd4818; ROM2[7491]<=16'd0; ROM3[7491]<=16'd23732; ROM4[7491]<=16'd57250;
ROM1[7492]<=16'd4810; ROM2[7492]<=16'd0; ROM3[7492]<=16'd23745; ROM4[7492]<=16'd57260;
ROM1[7493]<=16'd4816; ROM2[7493]<=16'd0; ROM3[7493]<=16'd23770; ROM4[7493]<=16'd57280;
ROM1[7494]<=16'd4808; ROM2[7494]<=16'd0; ROM3[7494]<=16'd23779; ROM4[7494]<=16'd57282;
ROM1[7495]<=16'd4787; ROM2[7495]<=16'd0; ROM3[7495]<=16'd23775; ROM4[7495]<=16'd57269;
ROM1[7496]<=16'd4772; ROM2[7496]<=16'd0; ROM3[7496]<=16'd23758; ROM4[7496]<=16'd57254;
ROM1[7497]<=16'd4781; ROM2[7497]<=16'd0; ROM3[7497]<=16'd23740; ROM4[7497]<=16'd57241;
ROM1[7498]<=16'd4810; ROM2[7498]<=16'd0; ROM3[7498]<=16'd23725; ROM4[7498]<=16'd57237;
ROM1[7499]<=16'd4820; ROM2[7499]<=16'd0; ROM3[7499]<=16'd23723; ROM4[7499]<=16'd57238;
ROM1[7500]<=16'd4821; ROM2[7500]<=16'd0; ROM3[7500]<=16'd23739; ROM4[7500]<=16'd57251;
ROM1[7501]<=16'd4816; ROM2[7501]<=16'd0; ROM3[7501]<=16'd23758; ROM4[7501]<=16'd57263;
ROM1[7502]<=16'd4798; ROM2[7502]<=16'd0; ROM3[7502]<=16'd23763; ROM4[7502]<=16'd57261;
ROM1[7503]<=16'd4780; ROM2[7503]<=16'd0; ROM3[7503]<=16'd23768; ROM4[7503]<=16'd57260;
ROM1[7504]<=16'd4769; ROM2[7504]<=16'd0; ROM3[7504]<=16'd23767; ROM4[7504]<=16'd57257;
ROM1[7505]<=16'd4785; ROM2[7505]<=16'd0; ROM3[7505]<=16'd23761; ROM4[7505]<=16'd57257;
ROM1[7506]<=16'd4822; ROM2[7506]<=16'd0; ROM3[7506]<=16'd23753; ROM4[7506]<=16'd57263;
ROM1[7507]<=16'd4850; ROM2[7507]<=16'd0; ROM3[7507]<=16'd23759; ROM4[7507]<=16'd57282;
ROM1[7508]<=16'd4840; ROM2[7508]<=16'd0; ROM3[7508]<=16'd23763; ROM4[7508]<=16'd57284;
ROM1[7509]<=16'd4804; ROM2[7509]<=16'd0; ROM3[7509]<=16'd23758; ROM4[7509]<=16'd57266;
ROM1[7510]<=16'd4792; ROM2[7510]<=16'd0; ROM3[7510]<=16'd23769; ROM4[7510]<=16'd57273;
ROM1[7511]<=16'd4781; ROM2[7511]<=16'd0; ROM3[7511]<=16'd23775; ROM4[7511]<=16'd57277;
ROM1[7512]<=16'd4767; ROM2[7512]<=16'd0; ROM3[7512]<=16'd23773; ROM4[7512]<=16'd57271;
ROM1[7513]<=16'd4777; ROM2[7513]<=16'd0; ROM3[7513]<=16'd23768; ROM4[7513]<=16'd57272;
ROM1[7514]<=16'd4815; ROM2[7514]<=16'd0; ROM3[7514]<=16'd23768; ROM4[7514]<=16'd57281;
ROM1[7515]<=16'd4840; ROM2[7515]<=16'd0; ROM3[7515]<=16'd23756; ROM4[7515]<=16'd57275;
ROM1[7516]<=16'd4831; ROM2[7516]<=16'd0; ROM3[7516]<=16'd23749; ROM4[7516]<=16'd57267;
ROM1[7517]<=16'd4819; ROM2[7517]<=16'd0; ROM3[7517]<=16'd23761; ROM4[7517]<=16'd57271;
ROM1[7518]<=16'd4798; ROM2[7518]<=16'd0; ROM3[7518]<=16'd23759; ROM4[7518]<=16'd57261;
ROM1[7519]<=16'd4795; ROM2[7519]<=16'd0; ROM3[7519]<=16'd23772; ROM4[7519]<=16'd57272;
ROM1[7520]<=16'd4787; ROM2[7520]<=16'd0; ROM3[7520]<=16'd23781; ROM4[7520]<=16'd57276;
ROM1[7521]<=16'd4771; ROM2[7521]<=16'd0; ROM3[7521]<=16'd23760; ROM4[7521]<=16'd57255;
ROM1[7522]<=16'd4787; ROM2[7522]<=16'd0; ROM3[7522]<=16'd23749; ROM4[7522]<=16'd57251;
ROM1[7523]<=16'd4813; ROM2[7523]<=16'd0; ROM3[7523]<=16'd23731; ROM4[7523]<=16'd57245;
ROM1[7524]<=16'd4824; ROM2[7524]<=16'd0; ROM3[7524]<=16'd23731; ROM4[7524]<=16'd57250;
ROM1[7525]<=16'd4833; ROM2[7525]<=16'd0; ROM3[7525]<=16'd23759; ROM4[7525]<=16'd57278;
ROM1[7526]<=16'd4818; ROM2[7526]<=16'd0; ROM3[7526]<=16'd23769; ROM4[7526]<=16'd57283;
ROM1[7527]<=16'd4792; ROM2[7527]<=16'd0; ROM3[7527]<=16'd23764; ROM4[7527]<=16'd57269;
ROM1[7528]<=16'd4774; ROM2[7528]<=16'd0; ROM3[7528]<=16'd23768; ROM4[7528]<=16'd57268;
ROM1[7529]<=16'd4776; ROM2[7529]<=16'd0; ROM3[7529]<=16'd23776; ROM4[7529]<=16'd57273;
ROM1[7530]<=16'd4795; ROM2[7530]<=16'd0; ROM3[7530]<=16'd23776; ROM4[7530]<=16'd57277;
ROM1[7531]<=16'd4820; ROM2[7531]<=16'd0; ROM3[7531]<=16'd23760; ROM4[7531]<=16'd57274;
ROM1[7532]<=16'd4837; ROM2[7532]<=16'd0; ROM3[7532]<=16'd23752; ROM4[7532]<=16'd57270;
ROM1[7533]<=16'd4834; ROM2[7533]<=16'd0; ROM3[7533]<=16'd23762; ROM4[7533]<=16'd57276;
ROM1[7534]<=16'd4821; ROM2[7534]<=16'd0; ROM3[7534]<=16'd23772; ROM4[7534]<=16'd57282;
ROM1[7535]<=16'd4805; ROM2[7535]<=16'd0; ROM3[7535]<=16'd23774; ROM4[7535]<=16'd57279;
ROM1[7536]<=16'd4800; ROM2[7536]<=16'd0; ROM3[7536]<=16'd23788; ROM4[7536]<=16'd57289;
ROM1[7537]<=16'd4817; ROM2[7537]<=16'd0; ROM3[7537]<=16'd23811; ROM4[7537]<=16'd57308;
ROM1[7538]<=16'd4821; ROM2[7538]<=16'd0; ROM3[7538]<=16'd23800; ROM4[7538]<=16'd57297;
ROM1[7539]<=16'd4833; ROM2[7539]<=16'd0; ROM3[7539]<=16'd23779; ROM4[7539]<=16'd57283;
ROM1[7540]<=16'd4847; ROM2[7540]<=16'd0; ROM3[7540]<=16'd23755; ROM4[7540]<=16'd57270;
ROM1[7541]<=16'd4833; ROM2[7541]<=16'd0; ROM3[7541]<=16'd23742; ROM4[7541]<=16'd57257;
ROM1[7542]<=16'd4832; ROM2[7542]<=16'd0; ROM3[7542]<=16'd23764; ROM4[7542]<=16'd57272;
ROM1[7543]<=16'd4829; ROM2[7543]<=16'd0; ROM3[7543]<=16'd23780; ROM4[7543]<=16'd57283;
ROM1[7544]<=16'd4804; ROM2[7544]<=16'd0; ROM3[7544]<=16'd23777; ROM4[7544]<=16'd57270;
ROM1[7545]<=16'd4774; ROM2[7545]<=16'd0; ROM3[7545]<=16'd23768; ROM4[7545]<=16'd57255;
ROM1[7546]<=16'd4769; ROM2[7546]<=16'd0; ROM3[7546]<=16'd23756; ROM4[7546]<=16'd57247;
ROM1[7547]<=16'd4797; ROM2[7547]<=16'd0; ROM3[7547]<=16'd23755; ROM4[7547]<=16'd57258;
ROM1[7548]<=16'd4836; ROM2[7548]<=16'd0; ROM3[7548]<=16'd23755; ROM4[7548]<=16'd57267;
ROM1[7549]<=16'd4838; ROM2[7549]<=16'd0; ROM3[7549]<=16'd23747; ROM4[7549]<=16'd57258;
ROM1[7550]<=16'd4821; ROM2[7550]<=16'd0; ROM3[7550]<=16'd23747; ROM4[7550]<=16'd57249;
ROM1[7551]<=16'd4803; ROM2[7551]<=16'd0; ROM3[7551]<=16'd23753; ROM4[7551]<=16'd57245;
ROM1[7552]<=16'd4792; ROM2[7552]<=16'd0; ROM3[7552]<=16'd23760; ROM4[7552]<=16'd57250;
ROM1[7553]<=16'd4780; ROM2[7553]<=16'd0; ROM3[7553]<=16'd23764; ROM4[7553]<=16'd57255;
ROM1[7554]<=16'd4777; ROM2[7554]<=16'd0; ROM3[7554]<=16'd23768; ROM4[7554]<=16'd57259;
ROM1[7555]<=16'd4798; ROM2[7555]<=16'd0; ROM3[7555]<=16'd23766; ROM4[7555]<=16'd57258;
ROM1[7556]<=16'd4839; ROM2[7556]<=16'd0; ROM3[7556]<=16'd23761; ROM4[7556]<=16'd57264;
ROM1[7557]<=16'd4866; ROM2[7557]<=16'd0; ROM3[7557]<=16'd23764; ROM4[7557]<=16'd57277;
ROM1[7558]<=16'd4856; ROM2[7558]<=16'd0; ROM3[7558]<=16'd23764; ROM4[7558]<=16'd57278;
ROM1[7559]<=16'd4840; ROM2[7559]<=16'd0; ROM3[7559]<=16'd23771; ROM4[7559]<=16'd57275;
ROM1[7560]<=16'd4832; ROM2[7560]<=16'd0; ROM3[7560]<=16'd23786; ROM4[7560]<=16'd57287;
ROM1[7561]<=16'd4827; ROM2[7561]<=16'd0; ROM3[7561]<=16'd23806; ROM4[7561]<=16'd57299;
ROM1[7562]<=16'd4797; ROM2[7562]<=16'd0; ROM3[7562]<=16'd23787; ROM4[7562]<=16'd57272;
ROM1[7563]<=16'd4782; ROM2[7563]<=16'd0; ROM3[7563]<=16'd23755; ROM4[7563]<=16'd57248;
ROM1[7564]<=16'd4800; ROM2[7564]<=16'd0; ROM3[7564]<=16'd23736; ROM4[7564]<=16'd57233;
ROM1[7565]<=16'd4812; ROM2[7565]<=16'd0; ROM3[7565]<=16'd23709; ROM4[7565]<=16'd57219;
ROM1[7566]<=16'd4816; ROM2[7566]<=16'd0; ROM3[7566]<=16'd23720; ROM4[7566]<=16'd57234;
ROM1[7567]<=16'd4811; ROM2[7567]<=16'd0; ROM3[7567]<=16'd23741; ROM4[7567]<=16'd57248;
ROM1[7568]<=16'd4793; ROM2[7568]<=16'd0; ROM3[7568]<=16'd23749; ROM4[7568]<=16'd57251;
ROM1[7569]<=16'd4776; ROM2[7569]<=16'd0; ROM3[7569]<=16'd23750; ROM4[7569]<=16'd57247;
ROM1[7570]<=16'd4770; ROM2[7570]<=16'd0; ROM3[7570]<=16'd23755; ROM4[7570]<=16'd57251;
ROM1[7571]<=16'd4780; ROM2[7571]<=16'd0; ROM3[7571]<=16'd23761; ROM4[7571]<=16'd57259;
ROM1[7572]<=16'd4801; ROM2[7572]<=16'd0; ROM3[7572]<=16'd23754; ROM4[7572]<=16'd57259;
ROM1[7573]<=16'd4845; ROM2[7573]<=16'd0; ROM3[7573]<=16'd23755; ROM4[7573]<=16'd57271;
ROM1[7574]<=16'd4867; ROM2[7574]<=16'd0; ROM3[7574]<=16'd23767; ROM4[7574]<=16'd57281;
ROM1[7575]<=16'd4845; ROM2[7575]<=16'd0; ROM3[7575]<=16'd23764; ROM4[7575]<=16'd57274;
ROM1[7576]<=16'd4810; ROM2[7576]<=16'd0; ROM3[7576]<=16'd23754; ROM4[7576]<=16'd57264;
ROM1[7577]<=16'd4781; ROM2[7577]<=16'd0; ROM3[7577]<=16'd23748; ROM4[7577]<=16'd57251;
ROM1[7578]<=16'd4764; ROM2[7578]<=16'd0; ROM3[7578]<=16'd23755; ROM4[7578]<=16'd57250;
ROM1[7579]<=16'd4769; ROM2[7579]<=16'd0; ROM3[7579]<=16'd23764; ROM4[7579]<=16'd57257;
ROM1[7580]<=16'd4796; ROM2[7580]<=16'd0; ROM3[7580]<=16'd23765; ROM4[7580]<=16'd57260;
ROM1[7581]<=16'd4833; ROM2[7581]<=16'd0; ROM3[7581]<=16'd23761; ROM4[7581]<=16'd57267;
ROM1[7582]<=16'd4849; ROM2[7582]<=16'd0; ROM3[7582]<=16'd23756; ROM4[7582]<=16'd57272;
ROM1[7583]<=16'd4845; ROM2[7583]<=16'd0; ROM3[7583]<=16'd23767; ROM4[7583]<=16'd57276;
ROM1[7584]<=16'd4838; ROM2[7584]<=16'd0; ROM3[7584]<=16'd23786; ROM4[7584]<=16'd57284;
ROM1[7585]<=16'd4823; ROM2[7585]<=16'd0; ROM3[7585]<=16'd23787; ROM4[7585]<=16'd57282;
ROM1[7586]<=16'd4810; ROM2[7586]<=16'd0; ROM3[7586]<=16'd23792; ROM4[7586]<=16'd57280;
ROM1[7587]<=16'd4818; ROM2[7587]<=16'd0; ROM3[7587]<=16'd23809; ROM4[7587]<=16'd57295;
ROM1[7588]<=16'd4835; ROM2[7588]<=16'd0; ROM3[7588]<=16'd23810; ROM4[7588]<=16'd57302;
ROM1[7589]<=16'd4859; ROM2[7589]<=16'd0; ROM3[7589]<=16'd23794; ROM4[7589]<=16'd57293;
ROM1[7590]<=16'd4890; ROM2[7590]<=16'd0; ROM3[7590]<=16'd23787; ROM4[7590]<=16'd57298;
ROM1[7591]<=16'd4889; ROM2[7591]<=16'd0; ROM3[7591]<=16'd23788; ROM4[7591]<=16'd57298;
ROM1[7592]<=16'd4871; ROM2[7592]<=16'd0; ROM3[7592]<=16'd23786; ROM4[7592]<=16'd57293;
ROM1[7593]<=16'd4855; ROM2[7593]<=16'd0; ROM3[7593]<=16'd23796; ROM4[7593]<=16'd57298;
ROM1[7594]<=16'd4837; ROM2[7594]<=16'd0; ROM3[7594]<=16'd23800; ROM4[7594]<=16'd57296;
ROM1[7595]<=16'd4814; ROM2[7595]<=16'd0; ROM3[7595]<=16'd23796; ROM4[7595]<=16'd57286;
ROM1[7596]<=16'd4813; ROM2[7596]<=16'd0; ROM3[7596]<=16'd23794; ROM4[7596]<=16'd57285;
ROM1[7597]<=16'd4839; ROM2[7597]<=16'd0; ROM3[7597]<=16'd23784; ROM4[7597]<=16'd57285;
ROM1[7598]<=16'd4870; ROM2[7598]<=16'd0; ROM3[7598]<=16'd23772; ROM4[7598]<=16'd57281;
ROM1[7599]<=16'd4879; ROM2[7599]<=16'd0; ROM3[7599]<=16'd23769; ROM4[7599]<=16'd57286;
ROM1[7600]<=16'd4874; ROM2[7600]<=16'd0; ROM3[7600]<=16'd23788; ROM4[7600]<=16'd57298;
ROM1[7601]<=16'd4867; ROM2[7601]<=16'd0; ROM3[7601]<=16'd23805; ROM4[7601]<=16'd57304;
ROM1[7602]<=16'd4857; ROM2[7602]<=16'd0; ROM3[7602]<=16'd23810; ROM4[7602]<=16'd57306;
ROM1[7603]<=16'd4832; ROM2[7603]<=16'd0; ROM3[7603]<=16'd23803; ROM4[7603]<=16'd57293;
ROM1[7604]<=16'd4841; ROM2[7604]<=16'd0; ROM3[7604]<=16'd23811; ROM4[7604]<=16'd57298;
ROM1[7605]<=16'd4870; ROM2[7605]<=16'd0; ROM3[7605]<=16'd23817; ROM4[7605]<=16'd57312;
ROM1[7606]<=16'd4882; ROM2[7606]<=16'd0; ROM3[7606]<=16'd23784; ROM4[7606]<=16'd57287;
ROM1[7607]<=16'd4880; ROM2[7607]<=16'd0; ROM3[7607]<=16'd23761; ROM4[7607]<=16'd57269;
ROM1[7608]<=16'd4858; ROM2[7608]<=16'd0; ROM3[7608]<=16'd23756; ROM4[7608]<=16'd57264;
ROM1[7609]<=16'd4823; ROM2[7609]<=16'd0; ROM3[7609]<=16'd23747; ROM4[7609]<=16'd57245;
ROM1[7610]<=16'd4812; ROM2[7610]<=16'd0; ROM3[7610]<=16'd23752; ROM4[7610]<=16'd57248;
ROM1[7611]<=16'd4810; ROM2[7611]<=16'd0; ROM3[7611]<=16'd23768; ROM4[7611]<=16'd57263;
ROM1[7612]<=16'd4801; ROM2[7612]<=16'd0; ROM3[7612]<=16'd23765; ROM4[7612]<=16'd57259;
ROM1[7613]<=16'd4805; ROM2[7613]<=16'd0; ROM3[7613]<=16'd23755; ROM4[7613]<=16'd57253;
ROM1[7614]<=16'd4831; ROM2[7614]<=16'd0; ROM3[7614]<=16'd23748; ROM4[7614]<=16'd57251;
ROM1[7615]<=16'd4855; ROM2[7615]<=16'd0; ROM3[7615]<=16'd23738; ROM4[7615]<=16'd57249;
ROM1[7616]<=16'd4851; ROM2[7616]<=16'd0; ROM3[7616]<=16'd23740; ROM4[7616]<=16'd57253;
ROM1[7617]<=16'd4830; ROM2[7617]<=16'd0; ROM3[7617]<=16'd23744; ROM4[7617]<=16'd57254;
ROM1[7618]<=16'd4820; ROM2[7618]<=16'd0; ROM3[7618]<=16'd23762; ROM4[7618]<=16'd57264;
ROM1[7619]<=16'd4827; ROM2[7619]<=16'd0; ROM3[7619]<=16'd23790; ROM4[7619]<=16'd57288;
ROM1[7620]<=16'd4807; ROM2[7620]<=16'd0; ROM3[7620]<=16'd23793; ROM4[7620]<=16'd57281;
ROM1[7621]<=16'd4797; ROM2[7621]<=16'd0; ROM3[7621]<=16'd23782; ROM4[7621]<=16'd57267;
ROM1[7622]<=16'd4818; ROM2[7622]<=16'd0; ROM3[7622]<=16'd23778; ROM4[7622]<=16'd57268;
ROM1[7623]<=16'd4847; ROM2[7623]<=16'd0; ROM3[7623]<=16'd23765; ROM4[7623]<=16'd57268;
ROM1[7624]<=16'd4847; ROM2[7624]<=16'd0; ROM3[7624]<=16'd23758; ROM4[7624]<=16'd57262;
ROM1[7625]<=16'd4840; ROM2[7625]<=16'd0; ROM3[7625]<=16'd23773; ROM4[7625]<=16'd57270;
ROM1[7626]<=16'd4840; ROM2[7626]<=16'd0; ROM3[7626]<=16'd23791; ROM4[7626]<=16'd57285;
ROM1[7627]<=16'd4834; ROM2[7627]<=16'd0; ROM3[7627]<=16'd23795; ROM4[7627]<=16'd57287;
ROM1[7628]<=16'd4799; ROM2[7628]<=16'd0; ROM3[7628]<=16'd23781; ROM4[7628]<=16'd57271;
ROM1[7629]<=16'd4784; ROM2[7629]<=16'd0; ROM3[7629]<=16'd23768; ROM4[7629]<=16'd57262;
ROM1[7630]<=16'd4805; ROM2[7630]<=16'd0; ROM3[7630]<=16'd23761; ROM4[7630]<=16'd57266;
ROM1[7631]<=16'd4842; ROM2[7631]<=16'd0; ROM3[7631]<=16'd23754; ROM4[7631]<=16'd57272;
ROM1[7632]<=16'd4882; ROM2[7632]<=16'd0; ROM3[7632]<=16'd23765; ROM4[7632]<=16'd57291;
ROM1[7633]<=16'd4887; ROM2[7633]<=16'd0; ROM3[7633]<=16'd23776; ROM4[7633]<=16'd57303;
ROM1[7634]<=16'd4855; ROM2[7634]<=16'd0; ROM3[7634]<=16'd23777; ROM4[7634]<=16'd57297;
ROM1[7635]<=16'd4833; ROM2[7635]<=16'd0; ROM3[7635]<=16'd23778; ROM4[7635]<=16'd57287;
ROM1[7636]<=16'd4829; ROM2[7636]<=16'd0; ROM3[7636]<=16'd23783; ROM4[7636]<=16'd57291;
ROM1[7637]<=16'd4825; ROM2[7637]<=16'd0; ROM3[7637]<=16'd23788; ROM4[7637]<=16'd57297;
ROM1[7638]<=16'd4848; ROM2[7638]<=16'd0; ROM3[7638]<=16'd23785; ROM4[7638]<=16'd57298;
ROM1[7639]<=16'd4897; ROM2[7639]<=16'd0; ROM3[7639]<=16'd23786; ROM4[7639]<=16'd57312;
ROM1[7640]<=16'd4928; ROM2[7640]<=16'd0; ROM3[7640]<=16'd23793; ROM4[7640]<=16'd57324;
ROM1[7641]<=16'd4915; ROM2[7641]<=16'd0; ROM3[7641]<=16'd23798; ROM4[7641]<=16'd57323;
ROM1[7642]<=16'd4900; ROM2[7642]<=16'd0; ROM3[7642]<=16'd23807; ROM4[7642]<=16'd57327;
ROM1[7643]<=16'd4873; ROM2[7643]<=16'd0; ROM3[7643]<=16'd23798; ROM4[7643]<=16'd57312;
ROM1[7644]<=16'd4866; ROM2[7644]<=16'd0; ROM3[7644]<=16'd23797; ROM4[7644]<=16'd57308;
ROM1[7645]<=16'd4860; ROM2[7645]<=16'd0; ROM3[7645]<=16'd23806; ROM4[7645]<=16'd57308;
ROM1[7646]<=16'd4857; ROM2[7646]<=16'd0; ROM3[7646]<=16'd23809; ROM4[7646]<=16'd57307;
ROM1[7647]<=16'd4930; ROM2[7647]<=16'd0; ROM3[7647]<=16'd23828; ROM4[7647]<=16'd57337;
ROM1[7648]<=16'd4971; ROM2[7648]<=16'd0; ROM3[7648]<=16'd23819; ROM4[7648]<=16'd57341;
ROM1[7649]<=16'd4988; ROM2[7649]<=16'd0; ROM3[7649]<=16'd23810; ROM4[7649]<=16'd57341;
ROM1[7650]<=16'd4994; ROM2[7650]<=16'd0; ROM3[7650]<=16'd23819; ROM4[7650]<=16'd57346;
ROM1[7651]<=16'd4962; ROM2[7651]<=16'd0; ROM3[7651]<=16'd23820; ROM4[7651]<=16'd57335;
ROM1[7652]<=16'd4971; ROM2[7652]<=16'd0; ROM3[7652]<=16'd23834; ROM4[7652]<=16'd57346;
ROM1[7653]<=16'd4992; ROM2[7653]<=16'd0; ROM3[7653]<=16'd23855; ROM4[7653]<=16'd57363;
ROM1[7654]<=16'd5019; ROM2[7654]<=16'd0; ROM3[7654]<=16'd23856; ROM4[7654]<=16'd57368;
ROM1[7655]<=16'd5053; ROM2[7655]<=16'd0; ROM3[7655]<=16'd23850; ROM4[7655]<=16'd57373;
ROM1[7656]<=16'd5106; ROM2[7656]<=16'd0; ROM3[7656]<=16'd23850; ROM4[7656]<=16'd57383;
ROM1[7657]<=16'd5149; ROM2[7657]<=16'd0; ROM3[7657]<=16'd23852; ROM4[7657]<=16'd57396;
ROM1[7658]<=16'd5172; ROM2[7658]<=16'd0; ROM3[7658]<=16'd23869; ROM4[7658]<=16'd57411;
ROM1[7659]<=16'd5167; ROM2[7659]<=16'd0; ROM3[7659]<=16'd23872; ROM4[7659]<=16'd57407;
ROM1[7660]<=16'd5175; ROM2[7660]<=16'd0; ROM3[7660]<=16'd23878; ROM4[7660]<=16'd57408;
ROM1[7661]<=16'd5215; ROM2[7661]<=16'd0; ROM3[7661]<=16'd23906; ROM4[7661]<=16'd57430;
ROM1[7662]<=16'd5222; ROM2[7662]<=16'd0; ROM3[7662]<=16'd23904; ROM4[7662]<=16'd57430;
ROM1[7663]<=16'd5225; ROM2[7663]<=16'd0; ROM3[7663]<=16'd23883; ROM4[7663]<=16'd57410;
ROM1[7664]<=16'd5257; ROM2[7664]<=16'd0; ROM3[7664]<=16'd23864; ROM4[7664]<=16'd57398;
ROM1[7665]<=16'd5288; ROM2[7665]<=16'd0; ROM3[7665]<=16'd23847; ROM4[7665]<=16'd57394;
ROM1[7666]<=16'd5300; ROM2[7666]<=16'd0; ROM3[7666]<=16'd23846; ROM4[7666]<=16'd57397;
ROM1[7667]<=16'd5319; ROM2[7667]<=16'd0; ROM3[7667]<=16'd23862; ROM4[7667]<=16'd57414;
ROM1[7668]<=16'd5321; ROM2[7668]<=16'd0; ROM3[7668]<=16'd23871; ROM4[7668]<=16'd57423;
ROM1[7669]<=16'd5307; ROM2[7669]<=16'd0; ROM3[7669]<=16'd23867; ROM4[7669]<=16'd57417;
ROM1[7670]<=16'd5299; ROM2[7670]<=16'd0; ROM3[7670]<=16'd23873; ROM4[7670]<=16'd57416;
ROM1[7671]<=16'd5314; ROM2[7671]<=16'd0; ROM3[7671]<=16'd23877; ROM4[7671]<=16'd57420;
ROM1[7672]<=16'd5350; ROM2[7672]<=16'd0; ROM3[7672]<=16'd23869; ROM4[7672]<=16'd57423;
ROM1[7673]<=16'd5398; ROM2[7673]<=16'd0; ROM3[7673]<=16'd23862; ROM4[7673]<=16'd57431;
ROM1[7674]<=16'd5434; ROM2[7674]<=16'd0; ROM3[7674]<=16'd23883; ROM4[7674]<=16'd57459;
ROM1[7675]<=16'd5454; ROM2[7675]<=16'd0; ROM3[7675]<=16'd23910; ROM4[7675]<=16'd57487;
ROM1[7676]<=16'd5439; ROM2[7676]<=16'd0; ROM3[7676]<=16'd23912; ROM4[7676]<=16'd57486;
ROM1[7677]<=16'd5436; ROM2[7677]<=16'd0; ROM3[7677]<=16'd23923; ROM4[7677]<=16'd57492;
ROM1[7678]<=16'd5436; ROM2[7678]<=16'd0; ROM3[7678]<=16'd23931; ROM4[7678]<=16'd57500;
ROM1[7679]<=16'd5417; ROM2[7679]<=16'd0; ROM3[7679]<=16'd23907; ROM4[7679]<=16'd57481;
ROM1[7680]<=16'd5438; ROM2[7680]<=16'd0; ROM3[7680]<=16'd23901; ROM4[7680]<=16'd57481;
ROM1[7681]<=16'd5469; ROM2[7681]<=16'd0; ROM3[7681]<=16'd23891; ROM4[7681]<=16'd57483;
ROM1[7682]<=16'd5480; ROM2[7682]<=16'd0; ROM3[7682]<=16'd23880; ROM4[7682]<=16'd57476;
ROM1[7683]<=16'd5480; ROM2[7683]<=16'd0; ROM3[7683]<=16'd23898; ROM4[7683]<=16'd57486;
ROM1[7684]<=16'd5487; ROM2[7684]<=16'd0; ROM3[7684]<=16'd23924; ROM4[7684]<=16'd57504;
ROM1[7685]<=16'd5475; ROM2[7685]<=16'd0; ROM3[7685]<=16'd23929; ROM4[7685]<=16'd57501;
ROM1[7686]<=16'd5443; ROM2[7686]<=16'd0; ROM3[7686]<=16'd23913; ROM4[7686]<=16'd57484;
ROM1[7687]<=16'd5431; ROM2[7687]<=16'd0; ROM3[7687]<=16'd23914; ROM4[7687]<=16'd57478;
ROM1[7688]<=16'd5440; ROM2[7688]<=16'd0; ROM3[7688]<=16'd23919; ROM4[7688]<=16'd57485;
ROM1[7689]<=16'd5464; ROM2[7689]<=16'd0; ROM3[7689]<=16'd23906; ROM4[7689]<=16'd57482;
ROM1[7690]<=16'd5494; ROM2[7690]<=16'd0; ROM3[7690]<=16'd23902; ROM4[7690]<=16'd57486;
ROM1[7691]<=16'd5491; ROM2[7691]<=16'd0; ROM3[7691]<=16'd23908; ROM4[7691]<=16'd57494;
ROM1[7692]<=16'd5462; ROM2[7692]<=16'd0; ROM3[7692]<=16'd23908; ROM4[7692]<=16'd57488;
ROM1[7693]<=16'd5442; ROM2[7693]<=16'd0; ROM3[7693]<=16'd23916; ROM4[7693]<=16'd57486;
ROM1[7694]<=16'd5423; ROM2[7694]<=16'd0; ROM3[7694]<=16'd23916; ROM4[7694]<=16'd57485;
ROM1[7695]<=16'd5406; ROM2[7695]<=16'd0; ROM3[7695]<=16'd23913; ROM4[7695]<=16'd57482;
ROM1[7696]<=16'd5398; ROM2[7696]<=16'd0; ROM3[7696]<=16'd23905; ROM4[7696]<=16'd57476;
ROM1[7697]<=16'd5412; ROM2[7697]<=16'd0; ROM3[7697]<=16'd23894; ROM4[7697]<=16'd57471;
ROM1[7698]<=16'd5437; ROM2[7698]<=16'd0; ROM3[7698]<=16'd23886; ROM4[7698]<=16'd57470;
ROM1[7699]<=16'd5435; ROM2[7699]<=16'd0; ROM3[7699]<=16'd23887; ROM4[7699]<=16'd57474;
ROM1[7700]<=16'd5428; ROM2[7700]<=16'd0; ROM3[7700]<=16'd23903; ROM4[7700]<=16'd57490;
ROM1[7701]<=16'd5397; ROM2[7701]<=16'd0; ROM3[7701]<=16'd23908; ROM4[7701]<=16'd57482;
ROM1[7702]<=16'd5361; ROM2[7702]<=16'd0; ROM3[7702]<=16'd23908; ROM4[7702]<=16'd57474;
ROM1[7703]<=16'd5325; ROM2[7703]<=16'd0; ROM3[7703]<=16'd23907; ROM4[7703]<=16'd57462;
ROM1[7704]<=16'd5294; ROM2[7704]<=16'd0; ROM3[7704]<=16'd23895; ROM4[7704]<=16'd57444;
ROM1[7705]<=16'd5302; ROM2[7705]<=16'd0; ROM3[7705]<=16'd23890; ROM4[7705]<=16'd57446;
ROM1[7706]<=16'd5325; ROM2[7706]<=16'd0; ROM3[7706]<=16'd23885; ROM4[7706]<=16'd57448;
ROM1[7707]<=16'd5316; ROM2[7707]<=16'd0; ROM3[7707]<=16'd23866; ROM4[7707]<=16'd57439;
ROM1[7708]<=16'd5283; ROM2[7708]<=16'd0; ROM3[7708]<=16'd23859; ROM4[7708]<=16'd57422;
ROM1[7709]<=16'd5255; ROM2[7709]<=16'd0; ROM3[7709]<=16'd23869; ROM4[7709]<=16'd57419;
ROM1[7710]<=16'd5230; ROM2[7710]<=16'd0; ROM3[7710]<=16'd23866; ROM4[7710]<=16'd57416;
ROM1[7711]<=16'd5215; ROM2[7711]<=16'd0; ROM3[7711]<=16'd23877; ROM4[7711]<=16'd57415;
ROM1[7712]<=16'd5218; ROM2[7712]<=16'd0; ROM3[7712]<=16'd23896; ROM4[7712]<=16'd57429;
ROM1[7713]<=16'd5233; ROM2[7713]<=16'd0; ROM3[7713]<=16'd23902; ROM4[7713]<=16'd57439;
ROM1[7714]<=16'd5248; ROM2[7714]<=16'd0; ROM3[7714]<=16'd23891; ROM4[7714]<=16'd57432;
ROM1[7715]<=16'd5247; ROM2[7715]<=16'd0; ROM3[7715]<=16'd23857; ROM4[7715]<=16'd57409;
ROM1[7716]<=16'd5217; ROM2[7716]<=16'd0; ROM3[7716]<=16'd23840; ROM4[7716]<=16'd57391;
ROM1[7717]<=16'd5175; ROM2[7717]<=16'd0; ROM3[7717]<=16'd23833; ROM4[7717]<=16'd57377;
ROM1[7718]<=16'd5148; ROM2[7718]<=16'd0; ROM3[7718]<=16'd23839; ROM4[7718]<=16'd57375;
ROM1[7719]<=16'd5132; ROM2[7719]<=16'd0; ROM3[7719]<=16'd23855; ROM4[7719]<=16'd57380;
ROM1[7720]<=16'd5101; ROM2[7720]<=16'd0; ROM3[7720]<=16'd23851; ROM4[7720]<=16'd57365;
ROM1[7721]<=16'd5091; ROM2[7721]<=16'd0; ROM3[7721]<=16'd23847; ROM4[7721]<=16'd57357;
ROM1[7722]<=16'd5111; ROM2[7722]<=16'd0; ROM3[7722]<=16'd23841; ROM4[7722]<=16'd57355;
ROM1[7723]<=16'd5148; ROM2[7723]<=16'd0; ROM3[7723]<=16'd23838; ROM4[7723]<=16'd57363;
ROM1[7724]<=16'd5147; ROM2[7724]<=16'd0; ROM3[7724]<=16'd23837; ROM4[7724]<=16'd57368;
ROM1[7725]<=16'd5124; ROM2[7725]<=16'd0; ROM3[7725]<=16'd23837; ROM4[7725]<=16'd57365;
ROM1[7726]<=16'd5108; ROM2[7726]<=16'd0; ROM3[7726]<=16'd23851; ROM4[7726]<=16'd57372;
ROM1[7727]<=16'd5087; ROM2[7727]<=16'd0; ROM3[7727]<=16'd23855; ROM4[7727]<=16'd57370;
ROM1[7728]<=16'd5055; ROM2[7728]<=16'd0; ROM3[7728]<=16'd23841; ROM4[7728]<=16'd57352;
ROM1[7729]<=16'd5039; ROM2[7729]<=16'd0; ROM3[7729]<=16'd23826; ROM4[7729]<=16'd57339;
ROM1[7730]<=16'd5044; ROM2[7730]<=16'd0; ROM3[7730]<=16'd23811; ROM4[7730]<=16'd57329;
ROM1[7731]<=16'd5076; ROM2[7731]<=16'd0; ROM3[7731]<=16'd23805; ROM4[7731]<=16'd57337;
ROM1[7732]<=16'd5112; ROM2[7732]<=16'd0; ROM3[7732]<=16'd23823; ROM4[7732]<=16'd57361;
ROM1[7733]<=16'd5095; ROM2[7733]<=16'd0; ROM3[7733]<=16'd23823; ROM4[7733]<=16'd57356;
ROM1[7734]<=16'd5062; ROM2[7734]<=16'd0; ROM3[7734]<=16'd23822; ROM4[7734]<=16'd57348;
ROM1[7735]<=16'd5043; ROM2[7735]<=16'd0; ROM3[7735]<=16'd23834; ROM4[7735]<=16'd57356;
ROM1[7736]<=16'd5026; ROM2[7736]<=16'd0; ROM3[7736]<=16'd23841; ROM4[7736]<=16'd57360;
ROM1[7737]<=16'd5026; ROM2[7737]<=16'd0; ROM3[7737]<=16'd23857; ROM4[7737]<=16'd57369;
ROM1[7738]<=16'd5037; ROM2[7738]<=16'd0; ROM3[7738]<=16'd23856; ROM4[7738]<=16'd57370;
ROM1[7739]<=16'd5073; ROM2[7739]<=16'd0; ROM3[7739]<=16'd23853; ROM4[7739]<=16'd57377;
ROM1[7740]<=16'd5107; ROM2[7740]<=16'd0; ROM3[7740]<=16'd23859; ROM4[7740]<=16'd57392;
ROM1[7741]<=16'd5091; ROM2[7741]<=16'd0; ROM3[7741]<=16'd23856; ROM4[7741]<=16'd57392;
ROM1[7742]<=16'd5056; ROM2[7742]<=16'd0; ROM3[7742]<=16'd23848; ROM4[7742]<=16'd57379;
ROM1[7743]<=16'd5026; ROM2[7743]<=16'd0; ROM3[7743]<=16'd23848; ROM4[7743]<=16'd57365;
ROM1[7744]<=16'd4998; ROM2[7744]<=16'd0; ROM3[7744]<=16'd23844; ROM4[7744]<=16'd57356;
ROM1[7745]<=16'd4984; ROM2[7745]<=16'd0; ROM3[7745]<=16'd23846; ROM4[7745]<=16'd57355;
ROM1[7746]<=16'd4999; ROM2[7746]<=16'd0; ROM3[7746]<=16'd23857; ROM4[7746]<=16'd57364;
ROM1[7747]<=16'd5025; ROM2[7747]<=16'd0; ROM3[7747]<=16'd23849; ROM4[7747]<=16'd57366;
ROM1[7748]<=16'd5061; ROM2[7748]<=16'd0; ROM3[7748]<=16'd23848; ROM4[7748]<=16'd57370;
ROM1[7749]<=16'd5058; ROM2[7749]<=16'd0; ROM3[7749]<=16'd23844; ROM4[7749]<=16'd57366;
ROM1[7750]<=16'd5028; ROM2[7750]<=16'd0; ROM3[7750]<=16'd23834; ROM4[7750]<=16'd57354;
ROM1[7751]<=16'd5012; ROM2[7751]<=16'd0; ROM3[7751]<=16'd23843; ROM4[7751]<=16'd57355;
ROM1[7752]<=16'd5003; ROM2[7752]<=16'd0; ROM3[7752]<=16'd23853; ROM4[7752]<=16'd57361;
ROM1[7753]<=16'd4989; ROM2[7753]<=16'd0; ROM3[7753]<=16'd23860; ROM4[7753]<=16'd57363;
ROM1[7754]<=16'd4986; ROM2[7754]<=16'd0; ROM3[7754]<=16'd23867; ROM4[7754]<=16'd57368;
ROM1[7755]<=16'd4999; ROM2[7755]<=16'd0; ROM3[7755]<=16'd23864; ROM4[7755]<=16'd57366;
ROM1[7756]<=16'd5028; ROM2[7756]<=16'd0; ROM3[7756]<=16'd23849; ROM4[7756]<=16'd57366;
ROM1[7757]<=16'd5056; ROM2[7757]<=16'd0; ROM3[7757]<=16'd23854; ROM4[7757]<=16'd57381;
ROM1[7758]<=16'd5052; ROM2[7758]<=16'd0; ROM3[7758]<=16'd23869; ROM4[7758]<=16'd57387;
ROM1[7759]<=16'd5008; ROM2[7759]<=16'd0; ROM3[7759]<=16'd23851; ROM4[7759]<=16'd57364;
ROM1[7760]<=16'd4964; ROM2[7760]<=16'd0; ROM3[7760]<=16'd23833; ROM4[7760]<=16'd57342;
ROM1[7761]<=16'd4935; ROM2[7761]<=16'd0; ROM3[7761]<=16'd23826; ROM4[7761]<=16'd57325;
ROM1[7762]<=16'd4927; ROM2[7762]<=16'd0; ROM3[7762]<=16'd23822; ROM4[7762]<=16'd57320;
ROM1[7763]<=16'd4947; ROM2[7763]<=16'd0; ROM3[7763]<=16'd23823; ROM4[7763]<=16'd57328;
ROM1[7764]<=16'd4975; ROM2[7764]<=16'd0; ROM3[7764]<=16'd23813; ROM4[7764]<=16'd57325;
ROM1[7765]<=16'd4993; ROM2[7765]<=16'd0; ROM3[7765]<=16'd23800; ROM4[7765]<=16'd57322;
ROM1[7766]<=16'd4982; ROM2[7766]<=16'd0; ROM3[7766]<=16'd23797; ROM4[7766]<=16'd57321;
ROM1[7767]<=16'd4963; ROM2[7767]<=16'd0; ROM3[7767]<=16'd23807; ROM4[7767]<=16'd57323;
ROM1[7768]<=16'd4943; ROM2[7768]<=16'd0; ROM3[7768]<=16'd23808; ROM4[7768]<=16'd57317;
ROM1[7769]<=16'd4929; ROM2[7769]<=16'd0; ROM3[7769]<=16'd23809; ROM4[7769]<=16'd57313;
ROM1[7770]<=16'd4913; ROM2[7770]<=16'd0; ROM3[7770]<=16'd23812; ROM4[7770]<=16'd57311;
ROM1[7771]<=16'd4905; ROM2[7771]<=16'd0; ROM3[7771]<=16'd23804; ROM4[7771]<=16'd57301;
ROM1[7772]<=16'd4936; ROM2[7772]<=16'd0; ROM3[7772]<=16'd23801; ROM4[7772]<=16'd57304;
ROM1[7773]<=16'd4977; ROM2[7773]<=16'd0; ROM3[7773]<=16'd23798; ROM4[7773]<=16'd57316;
ROM1[7774]<=16'd4963; ROM2[7774]<=16'd0; ROM3[7774]<=16'd23781; ROM4[7774]<=16'd57302;
ROM1[7775]<=16'd4932; ROM2[7775]<=16'd0; ROM3[7775]<=16'd23773; ROM4[7775]<=16'd57284;
ROM1[7776]<=16'd4917; ROM2[7776]<=16'd0; ROM3[7776]<=16'd23785; ROM4[7776]<=16'd57288;
ROM1[7777]<=16'd4907; ROM2[7777]<=16'd0; ROM3[7777]<=16'd23795; ROM4[7777]<=16'd57294;
ROM1[7778]<=16'd4897; ROM2[7778]<=16'd0; ROM3[7778]<=16'd23800; ROM4[7778]<=16'd57296;
ROM1[7779]<=16'd4899; ROM2[7779]<=16'd0; ROM3[7779]<=16'd23802; ROM4[7779]<=16'd57299;
ROM1[7780]<=16'd4921; ROM2[7780]<=16'd0; ROM3[7780]<=16'd23803; ROM4[7780]<=16'd57309;
ROM1[7781]<=16'd4950; ROM2[7781]<=16'd0; ROM3[7781]<=16'd23796; ROM4[7781]<=16'd57310;
ROM1[7782]<=16'd4979; ROM2[7782]<=16'd0; ROM3[7782]<=16'd23806; ROM4[7782]<=16'd57325;
ROM1[7783]<=16'd4985; ROM2[7783]<=16'd0; ROM3[7783]<=16'd23825; ROM4[7783]<=16'd57347;
ROM1[7784]<=16'd4943; ROM2[7784]<=16'd0; ROM3[7784]<=16'd23804; ROM4[7784]<=16'd57321;
ROM1[7785]<=16'd4906; ROM2[7785]<=16'd0; ROM3[7785]<=16'd23788; ROM4[7785]<=16'd57297;
ROM1[7786]<=16'd4886; ROM2[7786]<=16'd0; ROM3[7786]<=16'd23788; ROM4[7786]<=16'd57289;
ROM1[7787]<=16'd4872; ROM2[7787]<=16'd0; ROM3[7787]<=16'd23786; ROM4[7787]<=16'd57280;
ROM1[7788]<=16'd4884; ROM2[7788]<=16'd0; ROM3[7788]<=16'd23787; ROM4[7788]<=16'd57285;
ROM1[7789]<=16'd4924; ROM2[7789]<=16'd0; ROM3[7789]<=16'd23788; ROM4[7789]<=16'd57296;
ROM1[7790]<=16'd4958; ROM2[7790]<=16'd0; ROM3[7790]<=16'd23786; ROM4[7790]<=16'd57303;
ROM1[7791]<=16'd4946; ROM2[7791]<=16'd0; ROM3[7791]<=16'd23792; ROM4[7791]<=16'd57301;
ROM1[7792]<=16'd4920; ROM2[7792]<=16'd0; ROM3[7792]<=16'd23803; ROM4[7792]<=16'd57299;
ROM1[7793]<=16'd4900; ROM2[7793]<=16'd0; ROM3[7793]<=16'd23810; ROM4[7793]<=16'd57297;
ROM1[7794]<=16'd4893; ROM2[7794]<=16'd0; ROM3[7794]<=16'd23826; ROM4[7794]<=16'd57307;
ROM1[7795]<=16'd4895; ROM2[7795]<=16'd0; ROM3[7795]<=16'd23841; ROM4[7795]<=16'd57319;
ROM1[7796]<=16'd4904; ROM2[7796]<=16'd0; ROM3[7796]<=16'd23846; ROM4[7796]<=16'd57324;
ROM1[7797]<=16'd4923; ROM2[7797]<=16'd0; ROM3[7797]<=16'd23834; ROM4[7797]<=16'd57324;
ROM1[7798]<=16'd4948; ROM2[7798]<=16'd0; ROM3[7798]<=16'd23820; ROM4[7798]<=16'd57323;
ROM1[7799]<=16'd4947; ROM2[7799]<=16'd0; ROM3[7799]<=16'd23812; ROM4[7799]<=16'd57321;
ROM1[7800]<=16'd4943; ROM2[7800]<=16'd0; ROM3[7800]<=16'd23824; ROM4[7800]<=16'd57329;
ROM1[7801]<=16'd4938; ROM2[7801]<=16'd0; ROM3[7801]<=16'd23844; ROM4[7801]<=16'd57341;
ROM1[7802]<=16'd4935; ROM2[7802]<=16'd0; ROM3[7802]<=16'd23860; ROM4[7802]<=16'd57354;
ROM1[7803]<=16'd4907; ROM2[7803]<=16'd0; ROM3[7803]<=16'd23849; ROM4[7803]<=16'd57338;
ROM1[7804]<=16'd4893; ROM2[7804]<=16'd0; ROM3[7804]<=16'd23839; ROM4[7804]<=16'd57322;
ROM1[7805]<=16'd4928; ROM2[7805]<=16'd0; ROM3[7805]<=16'd23850; ROM4[7805]<=16'd57337;
ROM1[7806]<=16'd4940; ROM2[7806]<=16'd0; ROM3[7806]<=16'd23817; ROM4[7806]<=16'd57319;
ROM1[7807]<=16'd4949; ROM2[7807]<=16'd0; ROM3[7807]<=16'd23805; ROM4[7807]<=16'd57314;
ROM1[7808]<=16'd4943; ROM2[7808]<=16'd0; ROM3[7808]<=16'd23820; ROM4[7808]<=16'd57324;
ROM1[7809]<=16'd4918; ROM2[7809]<=16'd0; ROM3[7809]<=16'd23824; ROM4[7809]<=16'd57320;
ROM1[7810]<=16'd4891; ROM2[7810]<=16'd0; ROM3[7810]<=16'd23816; ROM4[7810]<=16'd57304;
ROM1[7811]<=16'd4873; ROM2[7811]<=16'd0; ROM3[7811]<=16'd23812; ROM4[7811]<=16'd57300;
ROM1[7812]<=16'd4870; ROM2[7812]<=16'd0; ROM3[7812]<=16'd23811; ROM4[7812]<=16'd57299;
ROM1[7813]<=16'd4870; ROM2[7813]<=16'd0; ROM3[7813]<=16'd23792; ROM4[7813]<=16'd57283;
ROM1[7814]<=16'd4903; ROM2[7814]<=16'd0; ROM3[7814]<=16'd23785; ROM4[7814]<=16'd57290;
ROM1[7815]<=16'd4937; ROM2[7815]<=16'd0; ROM3[7815]<=16'd23787; ROM4[7815]<=16'd57301;
ROM1[7816]<=16'd4920; ROM2[7816]<=16'd0; ROM3[7816]<=16'd23775; ROM4[7816]<=16'd57291;
ROM1[7817]<=16'd4895; ROM2[7817]<=16'd0; ROM3[7817]<=16'd23774; ROM4[7817]<=16'd57282;
ROM1[7818]<=16'd4897; ROM2[7818]<=16'd0; ROM3[7818]<=16'd23804; ROM4[7818]<=16'd57300;
ROM1[7819]<=16'd4887; ROM2[7819]<=16'd0; ROM3[7819]<=16'd23822; ROM4[7819]<=16'd57314;
ROM1[7820]<=16'd4865; ROM2[7820]<=16'd0; ROM3[7820]<=16'd23809; ROM4[7820]<=16'd57301;
ROM1[7821]<=16'd4859; ROM2[7821]<=16'd0; ROM3[7821]<=16'd23799; ROM4[7821]<=16'd57290;
ROM1[7822]<=16'd4877; ROM2[7822]<=16'd0; ROM3[7822]<=16'd23789; ROM4[7822]<=16'd57284;
ROM1[7823]<=16'd4915; ROM2[7823]<=16'd0; ROM3[7823]<=16'd23778; ROM4[7823]<=16'd57287;
ROM1[7824]<=16'd4934; ROM2[7824]<=16'd0; ROM3[7824]<=16'd23795; ROM4[7824]<=16'd57305;
ROM1[7825]<=16'd4923; ROM2[7825]<=16'd0; ROM3[7825]<=16'd23806; ROM4[7825]<=16'd57315;
ROM1[7826]<=16'd4903; ROM2[7826]<=16'd0; ROM3[7826]<=16'd23805; ROM4[7826]<=16'd57308;
ROM1[7827]<=16'd4886; ROM2[7827]<=16'd0; ROM3[7827]<=16'd23804; ROM4[7827]<=16'd57300;
ROM1[7828]<=16'd4888; ROM2[7828]<=16'd0; ROM3[7828]<=16'd23827; ROM4[7828]<=16'd57322;
ROM1[7829]<=16'd4908; ROM2[7829]<=16'd0; ROM3[7829]<=16'd23849; ROM4[7829]<=16'd57343;
ROM1[7830]<=16'd4888; ROM2[7830]<=16'd0; ROM3[7830]<=16'd23808; ROM4[7830]<=16'd57308;
ROM1[7831]<=16'd4889; ROM2[7831]<=16'd0; ROM3[7831]<=16'd23773; ROM4[7831]<=16'd57284;
ROM1[7832]<=16'd4896; ROM2[7832]<=16'd0; ROM3[7832]<=16'd23763; ROM4[7832]<=16'd57279;
ROM1[7833]<=16'd4876; ROM2[7833]<=16'd0; ROM3[7833]<=16'd23756; ROM4[7833]<=16'd57268;
ROM1[7834]<=16'd4872; ROM2[7834]<=16'd0; ROM3[7834]<=16'd23779; ROM4[7834]<=16'd57286;
ROM1[7835]<=16'd4871; ROM2[7835]<=16'd0; ROM3[7835]<=16'd23797; ROM4[7835]<=16'd57297;
ROM1[7836]<=16'd4843; ROM2[7836]<=16'd0; ROM3[7836]<=16'd23784; ROM4[7836]<=16'd57278;
ROM1[7837]<=16'd4824; ROM2[7837]<=16'd0; ROM3[7837]<=16'd23771; ROM4[7837]<=16'd57265;
ROM1[7838]<=16'd4849; ROM2[7838]<=16'd0; ROM3[7838]<=16'd23782; ROM4[7838]<=16'd57278;
ROM1[7839]<=16'd4888; ROM2[7839]<=16'd0; ROM3[7839]<=16'd23785; ROM4[7839]<=16'd57293;
ROM1[7840]<=16'd4910; ROM2[7840]<=16'd0; ROM3[7840]<=16'd23777; ROM4[7840]<=16'd57295;
ROM1[7841]<=16'd4900; ROM2[7841]<=16'd0; ROM3[7841]<=16'd23779; ROM4[7841]<=16'd57301;
ROM1[7842]<=16'd4892; ROM2[7842]<=16'd0; ROM3[7842]<=16'd23796; ROM4[7842]<=16'd57312;
ROM1[7843]<=16'd4880; ROM2[7843]<=16'd0; ROM3[7843]<=16'd23803; ROM4[7843]<=16'd57309;
ROM1[7844]<=16'd4848; ROM2[7844]<=16'd0; ROM3[7844]<=16'd23790; ROM4[7844]<=16'd57290;
ROM1[7845]<=16'd4819; ROM2[7845]<=16'd0; ROM3[7845]<=16'd23781; ROM4[7845]<=16'd57272;
ROM1[7846]<=16'd4822; ROM2[7846]<=16'd0; ROM3[7846]<=16'd23778; ROM4[7846]<=16'd57274;
ROM1[7847]<=16'd4847; ROM2[7847]<=16'd0; ROM3[7847]<=16'd23771; ROM4[7847]<=16'd57277;
ROM1[7848]<=16'd4882; ROM2[7848]<=16'd0; ROM3[7848]<=16'd23768; ROM4[7848]<=16'd57282;
ROM1[7849]<=16'd4902; ROM2[7849]<=16'd0; ROM3[7849]<=16'd23779; ROM4[7849]<=16'd57293;
ROM1[7850]<=16'd4894; ROM2[7850]<=16'd0; ROM3[7850]<=16'd23791; ROM4[7850]<=16'd57298;
ROM1[7851]<=16'd4874; ROM2[7851]<=16'd0; ROM3[7851]<=16'd23798; ROM4[7851]<=16'd57295;
ROM1[7852]<=16'd4854; ROM2[7852]<=16'd0; ROM3[7852]<=16'd23798; ROM4[7852]<=16'd57290;
ROM1[7853]<=16'd4843; ROM2[7853]<=16'd0; ROM3[7853]<=16'd23804; ROM4[7853]<=16'd57293;
ROM1[7854]<=16'd4844; ROM2[7854]<=16'd0; ROM3[7854]<=16'd23806; ROM4[7854]<=16'd57292;
ROM1[7855]<=16'd4863; ROM2[7855]<=16'd0; ROM3[7855]<=16'd23806; ROM4[7855]<=16'd57293;
ROM1[7856]<=16'd4899; ROM2[7856]<=16'd0; ROM3[7856]<=16'd23799; ROM4[7856]<=16'd57296;
ROM1[7857]<=16'd4904; ROM2[7857]<=16'd0; ROM3[7857]<=16'd23783; ROM4[7857]<=16'd57292;
ROM1[7858]<=16'd4883; ROM2[7858]<=16'd0; ROM3[7858]<=16'd23779; ROM4[7858]<=16'd57284;
ROM1[7859]<=16'd4861; ROM2[7859]<=16'd0; ROM3[7859]<=16'd23781; ROM4[7859]<=16'd57281;
ROM1[7860]<=16'd4852; ROM2[7860]<=16'd0; ROM3[7860]<=16'd23791; ROM4[7860]<=16'd57288;
ROM1[7861]<=16'd4841; ROM2[7861]<=16'd0; ROM3[7861]<=16'd23808; ROM4[7861]<=16'd57295;
ROM1[7862]<=16'd4826; ROM2[7862]<=16'd0; ROM3[7862]<=16'd23805; ROM4[7862]<=16'd57290;
ROM1[7863]<=16'd4823; ROM2[7863]<=16'd0; ROM3[7863]<=16'd23790; ROM4[7863]<=16'd57278;
ROM1[7864]<=16'd4854; ROM2[7864]<=16'd0; ROM3[7864]<=16'd23784; ROM4[7864]<=16'd57277;
ROM1[7865]<=16'd4873; ROM2[7865]<=16'd0; ROM3[7865]<=16'd23768; ROM4[7865]<=16'd57272;
ROM1[7866]<=16'd4853; ROM2[7866]<=16'd0; ROM3[7866]<=16'd23756; ROM4[7866]<=16'd57259;
ROM1[7867]<=16'd4841; ROM2[7867]<=16'd0; ROM3[7867]<=16'd23765; ROM4[7867]<=16'd57261;
ROM1[7868]<=16'd4843; ROM2[7868]<=16'd0; ROM3[7868]<=16'd23786; ROM4[7868]<=16'd57276;
ROM1[7869]<=16'd4837; ROM2[7869]<=16'd0; ROM3[7869]<=16'd23792; ROM4[7869]<=16'd57280;
ROM1[7870]<=16'd4820; ROM2[7870]<=16'd0; ROM3[7870]<=16'd23785; ROM4[7870]<=16'd57272;
ROM1[7871]<=16'd4825; ROM2[7871]<=16'd0; ROM3[7871]<=16'd23787; ROM4[7871]<=16'd57273;
ROM1[7872]<=16'd4839; ROM2[7872]<=16'd0; ROM3[7872]<=16'd23764; ROM4[7872]<=16'd57259;
ROM1[7873]<=16'd4864; ROM2[7873]<=16'd0; ROM3[7873]<=16'd23744; ROM4[7873]<=16'd57253;
ROM1[7874]<=16'd4868; ROM2[7874]<=16'd0; ROM3[7874]<=16'd23745; ROM4[7874]<=16'd57257;
ROM1[7875]<=16'd4850; ROM2[7875]<=16'd0; ROM3[7875]<=16'd23748; ROM4[7875]<=16'd57255;
ROM1[7876]<=16'd4823; ROM2[7876]<=16'd0; ROM3[7876]<=16'd23750; ROM4[7876]<=16'd57253;
ROM1[7877]<=16'd4812; ROM2[7877]<=16'd0; ROM3[7877]<=16'd23758; ROM4[7877]<=16'd57254;
ROM1[7878]<=16'd4808; ROM2[7878]<=16'd0; ROM3[7878]<=16'd23769; ROM4[7878]<=16'd57260;
ROM1[7879]<=16'd4811; ROM2[7879]<=16'd0; ROM3[7879]<=16'd23772; ROM4[7879]<=16'd57265;
ROM1[7880]<=16'd4831; ROM2[7880]<=16'd0; ROM3[7880]<=16'd23770; ROM4[7880]<=16'd57270;
ROM1[7881]<=16'd4856; ROM2[7881]<=16'd0; ROM3[7881]<=16'd23761; ROM4[7881]<=16'd57269;
ROM1[7882]<=16'd4864; ROM2[7882]<=16'd0; ROM3[7882]<=16'd23754; ROM4[7882]<=16'd57266;
ROM1[7883]<=16'd4857; ROM2[7883]<=16'd0; ROM3[7883]<=16'd23760; ROM4[7883]<=16'd57270;
ROM1[7884]<=16'd4846; ROM2[7884]<=16'd0; ROM3[7884]<=16'd23774; ROM4[7884]<=16'd57277;
ROM1[7885]<=16'd4856; ROM2[7885]<=16'd0; ROM3[7885]<=16'd23806; ROM4[7885]<=16'd57295;
ROM1[7886]<=16'd4843; ROM2[7886]<=16'd0; ROM3[7886]<=16'd23813; ROM4[7886]<=16'd57293;
ROM1[7887]<=16'd4794; ROM2[7887]<=16'd0; ROM3[7887]<=16'd23774; ROM4[7887]<=16'd57254;
ROM1[7888]<=16'd4804; ROM2[7888]<=16'd0; ROM3[7888]<=16'd23763; ROM4[7888]<=16'd57246;
ROM1[7889]<=16'd4834; ROM2[7889]<=16'd0; ROM3[7889]<=16'd23749; ROM4[7889]<=16'd57248;
ROM1[7890]<=16'd4845; ROM2[7890]<=16'd0; ROM3[7890]<=16'd23729; ROM4[7890]<=16'd57239;
ROM1[7891]<=16'd4850; ROM2[7891]<=16'd0; ROM3[7891]<=16'd23735; ROM4[7891]<=16'd57248;
ROM1[7892]<=16'd4832; ROM2[7892]<=16'd0; ROM3[7892]<=16'd23739; ROM4[7892]<=16'd57250;
ROM1[7893]<=16'd4804; ROM2[7893]<=16'd0; ROM3[7893]<=16'd23740; ROM4[7893]<=16'd57241;
ROM1[7894]<=16'd4801; ROM2[7894]<=16'd0; ROM3[7894]<=16'd23757; ROM4[7894]<=16'd57251;
ROM1[7895]<=16'd4814; ROM2[7895]<=16'd0; ROM3[7895]<=16'd23783; ROM4[7895]<=16'd57269;
ROM1[7896]<=16'd4821; ROM2[7896]<=16'd0; ROM3[7896]<=16'd23789; ROM4[7896]<=16'd57276;
ROM1[7897]<=16'd4829; ROM2[7897]<=16'd0; ROM3[7897]<=16'd23758; ROM4[7897]<=16'd57260;
ROM1[7898]<=16'd4842; ROM2[7898]<=16'd0; ROM3[7898]<=16'd23722; ROM4[7898]<=16'd57239;
ROM1[7899]<=16'd4846; ROM2[7899]<=16'd0; ROM3[7899]<=16'd23727; ROM4[7899]<=16'd57247;
ROM1[7900]<=16'd4825; ROM2[7900]<=16'd0; ROM3[7900]<=16'd23731; ROM4[7900]<=16'd57245;
ROM1[7901]<=16'd4802; ROM2[7901]<=16'd0; ROM3[7901]<=16'd23737; ROM4[7901]<=16'd57242;
ROM1[7902]<=16'd4802; ROM2[7902]<=16'd0; ROM3[7902]<=16'd23760; ROM4[7902]<=16'd57258;
ROM1[7903]<=16'd4791; ROM2[7903]<=16'd0; ROM3[7903]<=16'd23769; ROM4[7903]<=16'd57261;
ROM1[7904]<=16'd4785; ROM2[7904]<=16'd0; ROM3[7904]<=16'd23761; ROM4[7904]<=16'd57254;
ROM1[7905]<=16'd4813; ROM2[7905]<=16'd0; ROM3[7905]<=16'd23764; ROM4[7905]<=16'd57263;
ROM1[7906]<=16'd4849; ROM2[7906]<=16'd0; ROM3[7906]<=16'd23762; ROM4[7906]<=16'd57269;
ROM1[7907]<=16'd4855; ROM2[7907]<=16'd0; ROM3[7907]<=16'd23751; ROM4[7907]<=16'd57264;
ROM1[7908]<=16'd4851; ROM2[7908]<=16'd0; ROM3[7908]<=16'd23763; ROM4[7908]<=16'd57274;
ROM1[7909]<=16'd4845; ROM2[7909]<=16'd0; ROM3[7909]<=16'd23783; ROM4[7909]<=16'd57283;
ROM1[7910]<=16'd4837; ROM2[7910]<=16'd0; ROM3[7910]<=16'd23791; ROM4[7910]<=16'd57288;
ROM1[7911]<=16'd4828; ROM2[7911]<=16'd0; ROM3[7911]<=16'd23797; ROM4[7911]<=16'd57292;
ROM1[7912]<=16'd4819; ROM2[7912]<=16'd0; ROM3[7912]<=16'd23794; ROM4[7912]<=16'd57287;
ROM1[7913]<=16'd4822; ROM2[7913]<=16'd0; ROM3[7913]<=16'd23783; ROM4[7913]<=16'd57280;
ROM1[7914]<=16'd4857; ROM2[7914]<=16'd0; ROM3[7914]<=16'd23780; ROM4[7914]<=16'd57285;
ROM1[7915]<=16'd4902; ROM2[7915]<=16'd0; ROM3[7915]<=16'd23792; ROM4[7915]<=16'd57304;
ROM1[7916]<=16'd4897; ROM2[7916]<=16'd0; ROM3[7916]<=16'd23791; ROM4[7916]<=16'd57303;
ROM1[7917]<=16'd4868; ROM2[7917]<=16'd0; ROM3[7917]<=16'd23781; ROM4[7917]<=16'd57293;
ROM1[7918]<=16'd4842; ROM2[7918]<=16'd0; ROM3[7918]<=16'd23777; ROM4[7918]<=16'd57287;
ROM1[7919]<=16'd4816; ROM2[7919]<=16'd0; ROM3[7919]<=16'd23773; ROM4[7919]<=16'd57275;
ROM1[7920]<=16'd4814; ROM2[7920]<=16'd0; ROM3[7920]<=16'd23790; ROM4[7920]<=16'd57282;
ROM1[7921]<=16'd4817; ROM2[7921]<=16'd0; ROM3[7921]<=16'd23785; ROM4[7921]<=16'd57277;
ROM1[7922]<=16'd4837; ROM2[7922]<=16'd0; ROM3[7922]<=16'd23768; ROM4[7922]<=16'd57270;
ROM1[7923]<=16'd4867; ROM2[7923]<=16'd0; ROM3[7923]<=16'd23755; ROM4[7923]<=16'd57269;
ROM1[7924]<=16'd4863; ROM2[7924]<=16'd0; ROM3[7924]<=16'd23752; ROM4[7924]<=16'd57268;
ROM1[7925]<=16'd4859; ROM2[7925]<=16'd0; ROM3[7925]<=16'd23770; ROM4[7925]<=16'd57279;
ROM1[7926]<=16'd4853; ROM2[7926]<=16'd0; ROM3[7926]<=16'd23792; ROM4[7926]<=16'd57292;
ROM1[7927]<=16'd4843; ROM2[7927]<=16'd0; ROM3[7927]<=16'd23799; ROM4[7927]<=16'd57291;
ROM1[7928]<=16'd4823; ROM2[7928]<=16'd0; ROM3[7928]<=16'd23796; ROM4[7928]<=16'd57280;
ROM1[7929]<=16'd4818; ROM2[7929]<=16'd0; ROM3[7929]<=16'd23792; ROM4[7929]<=16'd57276;
ROM1[7930]<=16'd4845; ROM2[7930]<=16'd0; ROM3[7930]<=16'd23789; ROM4[7930]<=16'd57281;
ROM1[7931]<=16'd4875; ROM2[7931]<=16'd0; ROM3[7931]<=16'd23774; ROM4[7931]<=16'd57277;
ROM1[7932]<=16'd4878; ROM2[7932]<=16'd0; ROM3[7932]<=16'd23755; ROM4[7932]<=16'd57268;
ROM1[7933]<=16'd4875; ROM2[7933]<=16'd0; ROM3[7933]<=16'd23763; ROM4[7933]<=16'd57275;
ROM1[7934]<=16'd4867; ROM2[7934]<=16'd0; ROM3[7934]<=16'd23777; ROM4[7934]<=16'd57282;
ROM1[7935]<=16'd4839; ROM2[7935]<=16'd0; ROM3[7935]<=16'd23773; ROM4[7935]<=16'd57272;
ROM1[7936]<=16'd4809; ROM2[7936]<=16'd0; ROM3[7936]<=16'd23765; ROM4[7936]<=16'd57259;
ROM1[7937]<=16'd4814; ROM2[7937]<=16'd0; ROM3[7937]<=16'd23775; ROM4[7937]<=16'd57268;
ROM1[7938]<=16'd4820; ROM2[7938]<=16'd0; ROM3[7938]<=16'd23771; ROM4[7938]<=16'd57265;
ROM1[7939]<=16'd4831; ROM2[7939]<=16'd0; ROM3[7939]<=16'd23745; ROM4[7939]<=16'd57250;
ROM1[7940]<=16'd4863; ROM2[7940]<=16'd0; ROM3[7940]<=16'd23743; ROM4[7940]<=16'd57254;
ROM1[7941]<=16'd4855; ROM2[7941]<=16'd0; ROM3[7941]<=16'd23748; ROM4[7941]<=16'd57256;
ROM1[7942]<=16'd4838; ROM2[7942]<=16'd0; ROM3[7942]<=16'd23751; ROM4[7942]<=16'd57253;
ROM1[7943]<=16'd4832; ROM2[7943]<=16'd0; ROM3[7943]<=16'd23767; ROM4[7943]<=16'd57259;
ROM1[7944]<=16'd4820; ROM2[7944]<=16'd0; ROM3[7944]<=16'd23776; ROM4[7944]<=16'd57266;
ROM1[7945]<=16'd4804; ROM2[7945]<=16'd0; ROM3[7945]<=16'd23773; ROM4[7945]<=16'd57254;
ROM1[7946]<=16'd4802; ROM2[7946]<=16'd0; ROM3[7946]<=16'd23766; ROM4[7946]<=16'd57244;
ROM1[7947]<=16'd4831; ROM2[7947]<=16'd0; ROM3[7947]<=16'd23761; ROM4[7947]<=16'd57249;
ROM1[7948]<=16'd4868; ROM2[7948]<=16'd0; ROM3[7948]<=16'd23756; ROM4[7948]<=16'd57254;
ROM1[7949]<=16'd4872; ROM2[7949]<=16'd0; ROM3[7949]<=16'd23749; ROM4[7949]<=16'd57255;
ROM1[7950]<=16'd4853; ROM2[7950]<=16'd0; ROM3[7950]<=16'd23751; ROM4[7950]<=16'd57256;
ROM1[7951]<=16'd4853; ROM2[7951]<=16'd0; ROM3[7951]<=16'd23774; ROM4[7951]<=16'd57274;
ROM1[7952]<=16'd4851; ROM2[7952]<=16'd0; ROM3[7952]<=16'd23790; ROM4[7952]<=16'd57287;
ROM1[7953]<=16'd4809; ROM2[7953]<=16'd0; ROM3[7953]<=16'd23771; ROM4[7953]<=16'd57265;
ROM1[7954]<=16'd4798; ROM2[7954]<=16'd0; ROM3[7954]<=16'd23763; ROM4[7954]<=16'd57256;
ROM1[7955]<=16'd4819; ROM2[7955]<=16'd0; ROM3[7955]<=16'd23759; ROM4[7955]<=16'd57256;
ROM1[7956]<=16'd4854; ROM2[7956]<=16'd0; ROM3[7956]<=16'd23744; ROM4[7956]<=16'd57255;
ROM1[7957]<=16'd4883; ROM2[7957]<=16'd0; ROM3[7957]<=16'd23752; ROM4[7957]<=16'd57270;
ROM1[7958]<=16'd4876; ROM2[7958]<=16'd0; ROM3[7958]<=16'd23764; ROM4[7958]<=16'd57282;
ROM1[7959]<=16'd4853; ROM2[7959]<=16'd0; ROM3[7959]<=16'd23765; ROM4[7959]<=16'd57279;
ROM1[7960]<=16'd4832; ROM2[7960]<=16'd0; ROM3[7960]<=16'd23767; ROM4[7960]<=16'd57273;
ROM1[7961]<=16'd4821; ROM2[7961]<=16'd0; ROM3[7961]<=16'd23780; ROM4[7961]<=16'd57277;
ROM1[7962]<=16'd4825; ROM2[7962]<=16'd0; ROM3[7962]<=16'd23787; ROM4[7962]<=16'd57283;
ROM1[7963]<=16'd4844; ROM2[7963]<=16'd0; ROM3[7963]<=16'd23783; ROM4[7963]<=16'd57290;
ROM1[7964]<=16'd4876; ROM2[7964]<=16'd0; ROM3[7964]<=16'd23776; ROM4[7964]<=16'd57293;
ROM1[7965]<=16'd4889; ROM2[7965]<=16'd0; ROM3[7965]<=16'd23755; ROM4[7965]<=16'd57282;
ROM1[7966]<=16'd4872; ROM2[7966]<=16'd0; ROM3[7966]<=16'd23749; ROM4[7966]<=16'd57272;
ROM1[7967]<=16'd4852; ROM2[7967]<=16'd0; ROM3[7967]<=16'd23762; ROM4[7967]<=16'd57273;
ROM1[7968]<=16'd4824; ROM2[7968]<=16'd0; ROM3[7968]<=16'd23762; ROM4[7968]<=16'd57268;
ROM1[7969]<=16'd4818; ROM2[7969]<=16'd0; ROM3[7969]<=16'd23775; ROM4[7969]<=16'd57276;
ROM1[7970]<=16'd4812; ROM2[7970]<=16'd0; ROM3[7970]<=16'd23783; ROM4[7970]<=16'd57278;
ROM1[7971]<=16'd4810; ROM2[7971]<=16'd0; ROM3[7971]<=16'd23772; ROM4[7971]<=16'd57270;
ROM1[7972]<=16'd4838; ROM2[7972]<=16'd0; ROM3[7972]<=16'd23767; ROM4[7972]<=16'd57271;
ROM1[7973]<=16'd4864; ROM2[7973]<=16'd0; ROM3[7973]<=16'd23754; ROM4[7973]<=16'd57274;
ROM1[7974]<=16'd4856; ROM2[7974]<=16'd0; ROM3[7974]<=16'd23742; ROM4[7974]<=16'd57268;
ROM1[7975]<=16'd4842; ROM2[7975]<=16'd0; ROM3[7975]<=16'd23749; ROM4[7975]<=16'd57269;
ROM1[7976]<=16'd4830; ROM2[7976]<=16'd0; ROM3[7976]<=16'd23763; ROM4[7976]<=16'd57276;
ROM1[7977]<=16'd4818; ROM2[7977]<=16'd0; ROM3[7977]<=16'd23764; ROM4[7977]<=16'd57271;
ROM1[7978]<=16'd4812; ROM2[7978]<=16'd0; ROM3[7978]<=16'd23778; ROM4[7978]<=16'd57280;
ROM1[7979]<=16'd4820; ROM2[7979]<=16'd0; ROM3[7979]<=16'd23789; ROM4[7979]<=16'd57289;
ROM1[7980]<=16'd4867; ROM2[7980]<=16'd0; ROM3[7980]<=16'd23806; ROM4[7980]<=16'd57313;
ROM1[7981]<=16'd4886; ROM2[7981]<=16'd0; ROM3[7981]<=16'd23787; ROM4[7981]<=16'd57299;
ROM1[7982]<=16'd4859; ROM2[7982]<=16'd0; ROM3[7982]<=16'd23740; ROM4[7982]<=16'd57259;
ROM1[7983]<=16'd4840; ROM2[7983]<=16'd0; ROM3[7983]<=16'd23737; ROM4[7983]<=16'd57253;
ROM1[7984]<=16'd4813; ROM2[7984]<=16'd0; ROM3[7984]<=16'd23738; ROM4[7984]<=16'd57243;
ROM1[7985]<=16'd4804; ROM2[7985]<=16'd0; ROM3[7985]<=16'd23746; ROM4[7985]<=16'd57248;
ROM1[7986]<=16'd4809; ROM2[7986]<=16'd0; ROM3[7986]<=16'd23769; ROM4[7986]<=16'd57273;
ROM1[7987]<=16'd4806; ROM2[7987]<=16'd0; ROM3[7987]<=16'd23774; ROM4[7987]<=16'd57275;
ROM1[7988]<=16'd4806; ROM2[7988]<=16'd0; ROM3[7988]<=16'd23757; ROM4[7988]<=16'd57261;
ROM1[7989]<=16'd4835; ROM2[7989]<=16'd0; ROM3[7989]<=16'd23748; ROM4[7989]<=16'd57259;
ROM1[7990]<=16'd4865; ROM2[7990]<=16'd0; ROM3[7990]<=16'd23747; ROM4[7990]<=16'd57267;
ROM1[7991]<=16'd4858; ROM2[7991]<=16'd0; ROM3[7991]<=16'd23754; ROM4[7991]<=16'd57272;
ROM1[7992]<=16'd4834; ROM2[7992]<=16'd0; ROM3[7992]<=16'd23760; ROM4[7992]<=16'd57271;
ROM1[7993]<=16'd4822; ROM2[7993]<=16'd0; ROM3[7993]<=16'd23772; ROM4[7993]<=16'd57274;
ROM1[7994]<=16'd4820; ROM2[7994]<=16'd0; ROM3[7994]<=16'd23788; ROM4[7994]<=16'd57283;
ROM1[7995]<=16'd4808; ROM2[7995]<=16'd0; ROM3[7995]<=16'd23788; ROM4[7995]<=16'd57279;
ROM1[7996]<=16'd4813; ROM2[7996]<=16'd0; ROM3[7996]<=16'd23787; ROM4[7996]<=16'd57280;
ROM1[7997]<=16'd4836; ROM2[7997]<=16'd0; ROM3[7997]<=16'd23773; ROM4[7997]<=16'd57282;
ROM1[7998]<=16'd4867; ROM2[7998]<=16'd0; ROM3[7998]<=16'd23761; ROM4[7998]<=16'd57276;
ROM1[7999]<=16'd4881; ROM2[7999]<=16'd0; ROM3[7999]<=16'd23773; ROM4[7999]<=16'd57285;
ROM1[8000]<=16'd4867; ROM2[8000]<=16'd0; ROM3[8000]<=16'd23781; ROM4[8000]<=16'd57289;
ROM1[8001]<=16'd4850; ROM2[8001]<=16'd0; ROM3[8001]<=16'd23786; ROM4[8001]<=16'd57285;
ROM1[8002]<=16'd4846; ROM2[8002]<=16'd0; ROM3[8002]<=16'd23797; ROM4[8002]<=16'd57291;
ROM1[8003]<=16'd4814; ROM2[8003]<=16'd0; ROM3[8003]<=16'd23781; ROM4[8003]<=16'd57275;
ROM1[8004]<=16'd4801; ROM2[8004]<=16'd0; ROM3[8004]<=16'd23761; ROM4[8004]<=16'd57263;
ROM1[8005]<=16'd4834; ROM2[8005]<=16'd0; ROM3[8005]<=16'd23766; ROM4[8005]<=16'd57271;
ROM1[8006]<=16'd4861; ROM2[8006]<=16'd0; ROM3[8006]<=16'd23749; ROM4[8006]<=16'd57266;
ROM1[8007]<=16'd4869; ROM2[8007]<=16'd0; ROM3[8007]<=16'd23737; ROM4[8007]<=16'd57262;
ROM1[8008]<=16'd4867; ROM2[8008]<=16'd0; ROM3[8008]<=16'd23754; ROM4[8008]<=16'd57274;
ROM1[8009]<=16'd4850; ROM2[8009]<=16'd0; ROM3[8009]<=16'd23766; ROM4[8009]<=16'd57279;
ROM1[8010]<=16'd4840; ROM2[8010]<=16'd0; ROM3[8010]<=16'd23775; ROM4[8010]<=16'd57281;
ROM1[8011]<=16'd4829; ROM2[8011]<=16'd0; ROM3[8011]<=16'd23785; ROM4[8011]<=16'd57287;
ROM1[8012]<=16'd4827; ROM2[8012]<=16'd0; ROM3[8012]<=16'd23791; ROM4[8012]<=16'd57288;
ROM1[8013]<=16'd4838; ROM2[8013]<=16'd0; ROM3[8013]<=16'd23788; ROM4[8013]<=16'd57288;
ROM1[8014]<=16'd4863; ROM2[8014]<=16'd0; ROM3[8014]<=16'd23781; ROM4[8014]<=16'd57290;
ROM1[8015]<=16'd4889; ROM2[8015]<=16'd0; ROM3[8015]<=16'd23772; ROM4[8015]<=16'd57292;
ROM1[8016]<=16'd4887; ROM2[8016]<=16'd0; ROM3[8016]<=16'd23774; ROM4[8016]<=16'd57293;
ROM1[8017]<=16'd4867; ROM2[8017]<=16'd0; ROM3[8017]<=16'd23782; ROM4[8017]<=16'd57296;
ROM1[8018]<=16'd4847; ROM2[8018]<=16'd0; ROM3[8018]<=16'd23791; ROM4[8018]<=16'd57298;
ROM1[8019]<=16'd4834; ROM2[8019]<=16'd0; ROM3[8019]<=16'd23801; ROM4[8019]<=16'd57300;
ROM1[8020]<=16'd4825; ROM2[8020]<=16'd0; ROM3[8020]<=16'd23810; ROM4[8020]<=16'd57304;
ROM1[8021]<=16'd4831; ROM2[8021]<=16'd0; ROM3[8021]<=16'd23807; ROM4[8021]<=16'd57305;
ROM1[8022]<=16'd4855; ROM2[8022]<=16'd0; ROM3[8022]<=16'd23798; ROM4[8022]<=16'd57301;
ROM1[8023]<=16'd4888; ROM2[8023]<=16'd0; ROM3[8023]<=16'd23791; ROM4[8023]<=16'd57303;
ROM1[8024]<=16'd4892; ROM2[8024]<=16'd0; ROM3[8024]<=16'd23793; ROM4[8024]<=16'd57311;
ROM1[8025]<=16'd4895; ROM2[8025]<=16'd0; ROM3[8025]<=16'd23819; ROM4[8025]<=16'd57329;
ROM1[8026]<=16'd4884; ROM2[8026]<=16'd0; ROM3[8026]<=16'd23832; ROM4[8026]<=16'd57336;
ROM1[8027]<=16'd4846; ROM2[8027]<=16'd0; ROM3[8027]<=16'd23819; ROM4[8027]<=16'd57318;
ROM1[8028]<=16'd4825; ROM2[8028]<=16'd0; ROM3[8028]<=16'd23816; ROM4[8028]<=16'd57311;
ROM1[8029]<=16'd4816; ROM2[8029]<=16'd0; ROM3[8029]<=16'd23809; ROM4[8029]<=16'd57304;
ROM1[8030]<=16'd4829; ROM2[8030]<=16'd0; ROM3[8030]<=16'd23797; ROM4[8030]<=16'd57297;
ROM1[8031]<=16'd4873; ROM2[8031]<=16'd0; ROM3[8031]<=16'd23791; ROM4[8031]<=16'd57307;
ROM1[8032]<=16'd4892; ROM2[8032]<=16'd0; ROM3[8032]<=16'd23795; ROM4[8032]<=16'd57313;
ROM1[8033]<=16'd4889; ROM2[8033]<=16'd0; ROM3[8033]<=16'd23811; ROM4[8033]<=16'd57326;
ROM1[8034]<=16'd4869; ROM2[8034]<=16'd0; ROM3[8034]<=16'd23817; ROM4[8034]<=16'd57329;
ROM1[8035]<=16'd4845; ROM2[8035]<=16'd0; ROM3[8035]<=16'd23811; ROM4[8035]<=16'd57317;
ROM1[8036]<=16'd4822; ROM2[8036]<=16'd0; ROM3[8036]<=16'd23805; ROM4[8036]<=16'd57305;
ROM1[8037]<=16'd4806; ROM2[8037]<=16'd0; ROM3[8037]<=16'd23794; ROM4[8037]<=16'd57288;
ROM1[8038]<=16'd4835; ROM2[8038]<=16'd0; ROM3[8038]<=16'd23798; ROM4[8038]<=16'd57299;
ROM1[8039]<=16'd4882; ROM2[8039]<=16'd0; ROM3[8039]<=16'd23797; ROM4[8039]<=16'd57312;
ROM1[8040]<=16'd4891; ROM2[8040]<=16'd0; ROM3[8040]<=16'd23771; ROM4[8040]<=16'd57297;
ROM1[8041]<=16'd4875; ROM2[8041]<=16'd0; ROM3[8041]<=16'd23760; ROM4[8041]<=16'd57285;
ROM1[8042]<=16'd4846; ROM2[8042]<=16'd0; ROM3[8042]<=16'd23759; ROM4[8042]<=16'd57273;
ROM1[8043]<=16'd4831; ROM2[8043]<=16'd0; ROM3[8043]<=16'd23766; ROM4[8043]<=16'd57274;
ROM1[8044]<=16'd4827; ROM2[8044]<=16'd0; ROM3[8044]<=16'd23778; ROM4[8044]<=16'd57285;
ROM1[8045]<=16'd4818; ROM2[8045]<=16'd0; ROM3[8045]<=16'd23784; ROM4[8045]<=16'd57287;
ROM1[8046]<=16'd4831; ROM2[8046]<=16'd0; ROM3[8046]<=16'd23782; ROM4[8046]<=16'd57287;
ROM1[8047]<=16'd4873; ROM2[8047]<=16'd0; ROM3[8047]<=16'd23786; ROM4[8047]<=16'd57299;
ROM1[8048]<=16'd4907; ROM2[8048]<=16'd0; ROM3[8048]<=16'd23781; ROM4[8048]<=16'd57302;
ROM1[8049]<=16'd4898; ROM2[8049]<=16'd0; ROM3[8049]<=16'd23770; ROM4[8049]<=16'd57291;
ROM1[8050]<=16'd4869; ROM2[8050]<=16'd0; ROM3[8050]<=16'd23768; ROM4[8050]<=16'd57283;
ROM1[8051]<=16'd4845; ROM2[8051]<=16'd0; ROM3[8051]<=16'd23775; ROM4[8051]<=16'd57279;
ROM1[8052]<=16'd4831; ROM2[8052]<=16'd0; ROM3[8052]<=16'd23784; ROM4[8052]<=16'd57283;
ROM1[8053]<=16'd4823; ROM2[8053]<=16'd0; ROM3[8053]<=16'd23799; ROM4[8053]<=16'd57292;
ROM1[8054]<=16'd4833; ROM2[8054]<=16'd0; ROM3[8054]<=16'd23808; ROM4[8054]<=16'd57302;
ROM1[8055]<=16'd4854; ROM2[8055]<=16'd0; ROM3[8055]<=16'd23803; ROM4[8055]<=16'd57300;
ROM1[8056]<=16'd4890; ROM2[8056]<=16'd0; ROM3[8056]<=16'd23799; ROM4[8056]<=16'd57301;
ROM1[8057]<=16'd4918; ROM2[8057]<=16'd0; ROM3[8057]<=16'd23804; ROM4[8057]<=16'd57316;
ROM1[8058]<=16'd4895; ROM2[8058]<=16'd0; ROM3[8058]<=16'd23804; ROM4[8058]<=16'd57310;
ROM1[8059]<=16'd4855; ROM2[8059]<=16'd0; ROM3[8059]<=16'd23797; ROM4[8059]<=16'd57297;
ROM1[8060]<=16'd4836; ROM2[8060]<=16'd0; ROM3[8060]<=16'd23795; ROM4[8060]<=16'd57295;
ROM1[8061]<=16'd4835; ROM2[8061]<=16'd0; ROM3[8061]<=16'd23811; ROM4[8061]<=16'd57307;
ROM1[8062]<=16'd4869; ROM2[8062]<=16'd0; ROM3[8062]<=16'd23845; ROM4[8062]<=16'd57345;
ROM1[8063]<=16'd4890; ROM2[8063]<=16'd0; ROM3[8063]<=16'd23852; ROM4[8063]<=16'd57355;
ROM1[8064]<=16'd4909; ROM2[8064]<=16'd0; ROM3[8064]<=16'd23829; ROM4[8064]<=16'd57340;
ROM1[8065]<=16'd4924; ROM2[8065]<=16'd0; ROM3[8065]<=16'd23810; ROM4[8065]<=16'd57332;
ROM1[8066]<=16'd4904; ROM2[8066]<=16'd0; ROM3[8066]<=16'd23800; ROM4[8066]<=16'd57321;
ROM1[8067]<=16'd4889; ROM2[8067]<=16'd0; ROM3[8067]<=16'd23810; ROM4[8067]<=16'd57324;
ROM1[8068]<=16'd4886; ROM2[8068]<=16'd0; ROM3[8068]<=16'd23837; ROM4[8068]<=16'd57341;
ROM1[8069]<=16'd4877; ROM2[8069]<=16'd0; ROM3[8069]<=16'd23851; ROM4[8069]<=16'd57347;
ROM1[8070]<=16'd4862; ROM2[8070]<=16'd0; ROM3[8070]<=16'd23851; ROM4[8070]<=16'd57342;
ROM1[8071]<=16'd4869; ROM2[8071]<=16'd0; ROM3[8071]<=16'd23854; ROM4[8071]<=16'd57345;
ROM1[8072]<=16'd4897; ROM2[8072]<=16'd0; ROM3[8072]<=16'd23848; ROM4[8072]<=16'd57349;
ROM1[8073]<=16'd4921; ROM2[8073]<=16'd0; ROM3[8073]<=16'd23828; ROM4[8073]<=16'd57346;
ROM1[8074]<=16'd4921; ROM2[8074]<=16'd0; ROM3[8074]<=16'd23820; ROM4[8074]<=16'd57338;
ROM1[8075]<=16'd4902; ROM2[8075]<=16'd0; ROM3[8075]<=16'd23824; ROM4[8075]<=16'd57335;
ROM1[8076]<=16'd4883; ROM2[8076]<=16'd0; ROM3[8076]<=16'd23829; ROM4[8076]<=16'd57334;
ROM1[8077]<=16'd4875; ROM2[8077]<=16'd0; ROM3[8077]<=16'd23840; ROM4[8077]<=16'd57341;
ROM1[8078]<=16'd4879; ROM2[8078]<=16'd0; ROM3[8078]<=16'd23857; ROM4[8078]<=16'd57361;
ROM1[8079]<=16'd4888; ROM2[8079]<=16'd0; ROM3[8079]<=16'd23857; ROM4[8079]<=16'd57367;
ROM1[8080]<=16'd4885; ROM2[8080]<=16'd0; ROM3[8080]<=16'd23828; ROM4[8080]<=16'd57345;
ROM1[8081]<=16'd4902; ROM2[8081]<=16'd0; ROM3[8081]<=16'd23806; ROM4[8081]<=16'd57334;
ROM1[8082]<=16'd4906; ROM2[8082]<=16'd0; ROM3[8082]<=16'd23794; ROM4[8082]<=16'd57327;
ROM1[8083]<=16'd4896; ROM2[8083]<=16'd0; ROM3[8083]<=16'd23796; ROM4[8083]<=16'd57331;
ROM1[8084]<=16'd4898; ROM2[8084]<=16'd0; ROM3[8084]<=16'd23822; ROM4[8084]<=16'd57350;
ROM1[8085]<=16'd4898; ROM2[8085]<=16'd0; ROM3[8085]<=16'd23844; ROM4[8085]<=16'd57360;
ROM1[8086]<=16'd4866; ROM2[8086]<=16'd0; ROM3[8086]<=16'd23838; ROM4[8086]<=16'd57349;
ROM1[8087]<=16'd4820; ROM2[8087]<=16'd0; ROM3[8087]<=16'd23801; ROM4[8087]<=16'd57309;
ROM1[8088]<=16'd4829; ROM2[8088]<=16'd0; ROM3[8088]<=16'd23784; ROM4[8088]<=16'd57295;
ROM1[8089]<=16'd4865; ROM2[8089]<=16'd0; ROM3[8089]<=16'd23775; ROM4[8089]<=16'd57300;
ROM1[8090]<=16'd4880; ROM2[8090]<=16'd0; ROM3[8090]<=16'd23758; ROM4[8090]<=16'd57291;
ROM1[8091]<=16'd4883; ROM2[8091]<=16'd0; ROM3[8091]<=16'd23769; ROM4[8091]<=16'd57298;
ROM1[8092]<=16'd4863; ROM2[8092]<=16'd0; ROM3[8092]<=16'd23779; ROM4[8092]<=16'd57303;
ROM1[8093]<=16'd4825; ROM2[8093]<=16'd0; ROM3[8093]<=16'd23772; ROM4[8093]<=16'd57287;
ROM1[8094]<=16'd4810; ROM2[8094]<=16'd0; ROM3[8094]<=16'd23778; ROM4[8094]<=16'd57284;
ROM1[8095]<=16'd4809; ROM2[8095]<=16'd0; ROM3[8095]<=16'd23788; ROM4[8095]<=16'd57288;
ROM1[8096]<=16'd4823; ROM2[8096]<=16'd0; ROM3[8096]<=16'd23796; ROM4[8096]<=16'd57300;
ROM1[8097]<=16'd4848; ROM2[8097]<=16'd0; ROM3[8097]<=16'd23784; ROM4[8097]<=16'd57296;
ROM1[8098]<=16'd4873; ROM2[8098]<=16'd0; ROM3[8098]<=16'd23765; ROM4[8098]<=16'd57288;
ROM1[8099]<=16'd4870; ROM2[8099]<=16'd0; ROM3[8099]<=16'd23758; ROM4[8099]<=16'd57286;
ROM1[8100]<=16'd4842; ROM2[8100]<=16'd0; ROM3[8100]<=16'd23751; ROM4[8100]<=16'd57272;
ROM1[8101]<=16'd4824; ROM2[8101]<=16'd0; ROM3[8101]<=16'd23761; ROM4[8101]<=16'd57272;
ROM1[8102]<=16'd4819; ROM2[8102]<=16'd0; ROM3[8102]<=16'd23770; ROM4[8102]<=16'd57281;
ROM1[8103]<=16'd4809; ROM2[8103]<=16'd0; ROM3[8103]<=16'd23779; ROM4[8103]<=16'd57285;
ROM1[8104]<=16'd4811; ROM2[8104]<=16'd0; ROM3[8104]<=16'd23780; ROM4[8104]<=16'd57286;
ROM1[8105]<=16'd4836; ROM2[8105]<=16'd0; ROM3[8105]<=16'd23780; ROM4[8105]<=16'd57289;
ROM1[8106]<=16'd4869; ROM2[8106]<=16'd0; ROM3[8106]<=16'd23769; ROM4[8106]<=16'd57290;
ROM1[8107]<=16'd4879; ROM2[8107]<=16'd0; ROM3[8107]<=16'd23763; ROM4[8107]<=16'd57291;
ROM1[8108]<=16'd4869; ROM2[8108]<=16'd0; ROM3[8108]<=16'd23768; ROM4[8108]<=16'd57294;
ROM1[8109]<=16'd4849; ROM2[8109]<=16'd0; ROM3[8109]<=16'd23772; ROM4[8109]<=16'd57294;
ROM1[8110]<=16'd4829; ROM2[8110]<=16'd0; ROM3[8110]<=16'd23779; ROM4[8110]<=16'd57292;
ROM1[8111]<=16'd4817; ROM2[8111]<=16'd0; ROM3[8111]<=16'd23790; ROM4[8111]<=16'd57295;
ROM1[8112]<=16'd4812; ROM2[8112]<=16'd0; ROM3[8112]<=16'd23791; ROM4[8112]<=16'd57295;
ROM1[8113]<=16'd4822; ROM2[8113]<=16'd0; ROM3[8113]<=16'd23784; ROM4[8113]<=16'd57289;
ROM1[8114]<=16'd4861; ROM2[8114]<=16'd0; ROM3[8114]<=16'd23785; ROM4[8114]<=16'd57296;
ROM1[8115]<=16'd4884; ROM2[8115]<=16'd0; ROM3[8115]<=16'd23780; ROM4[8115]<=16'd57296;
ROM1[8116]<=16'd4870; ROM2[8116]<=16'd0; ROM3[8116]<=16'd23776; ROM4[8116]<=16'd57288;
ROM1[8117]<=16'd4849; ROM2[8117]<=16'd0; ROM3[8117]<=16'd23782; ROM4[8117]<=16'd57286;
ROM1[8118]<=16'd4828; ROM2[8118]<=16'd0; ROM3[8118]<=16'd23784; ROM4[8118]<=16'd57285;
ROM1[8119]<=16'd4814; ROM2[8119]<=16'd0; ROM3[8119]<=16'd23786; ROM4[8119]<=16'd57285;
ROM1[8120]<=16'd4804; ROM2[8120]<=16'd0; ROM3[8120]<=16'd23795; ROM4[8120]<=16'd57290;
ROM1[8121]<=16'd4810; ROM2[8121]<=16'd0; ROM3[8121]<=16'd23795; ROM4[8121]<=16'd57292;
ROM1[8122]<=16'd4838; ROM2[8122]<=16'd0; ROM3[8122]<=16'd23785; ROM4[8122]<=16'd57294;
ROM1[8123]<=16'd4877; ROM2[8123]<=16'd0; ROM3[8123]<=16'd23782; ROM4[8123]<=16'd57305;
ROM1[8124]<=16'd4888; ROM2[8124]<=16'd0; ROM3[8124]<=16'd23789; ROM4[8124]<=16'd57312;
ROM1[8125]<=16'd4878; ROM2[8125]<=16'd0; ROM3[8125]<=16'd23802; ROM4[8125]<=16'd57322;
ROM1[8126]<=16'd4865; ROM2[8126]<=16'd0; ROM3[8126]<=16'd23817; ROM4[8126]<=16'd57329;
ROM1[8127]<=16'd4844; ROM2[8127]<=16'd0; ROM3[8127]<=16'd23817; ROM4[8127]<=16'd57320;
ROM1[8128]<=16'd4818; ROM2[8128]<=16'd0; ROM3[8128]<=16'd23810; ROM4[8128]<=16'd57311;
ROM1[8129]<=16'd4815; ROM2[8129]<=16'd0; ROM3[8129]<=16'd23804; ROM4[8129]<=16'd57307;
ROM1[8130]<=16'd4830; ROM2[8130]<=16'd0; ROM3[8130]<=16'd23796; ROM4[8130]<=16'd57302;
ROM1[8131]<=16'd4865; ROM2[8131]<=16'd0; ROM3[8131]<=16'd23785; ROM4[8131]<=16'd57308;
ROM1[8132]<=16'd4883; ROM2[8132]<=16'd0; ROM3[8132]<=16'd23786; ROM4[8132]<=16'd57314;
ROM1[8133]<=16'd4864; ROM2[8133]<=16'd0; ROM3[8133]<=16'd23783; ROM4[8133]<=16'd57304;
ROM1[8134]<=16'd4845; ROM2[8134]<=16'd0; ROM3[8134]<=16'd23791; ROM4[8134]<=16'd57297;
ROM1[8135]<=16'd4841; ROM2[8135]<=16'd0; ROM3[8135]<=16'd23805; ROM4[8135]<=16'd57302;
ROM1[8136]<=16'd4841; ROM2[8136]<=16'd0; ROM3[8136]<=16'd23820; ROM4[8136]<=16'd57316;
ROM1[8137]<=16'd4826; ROM2[8137]<=16'd0; ROM3[8137]<=16'd23812; ROM4[8137]<=16'd57305;
ROM1[8138]<=16'd4820; ROM2[8138]<=16'd0; ROM3[8138]<=16'd23786; ROM4[8138]<=16'd57285;
ROM1[8139]<=16'd4852; ROM2[8139]<=16'd0; ROM3[8139]<=16'd23775; ROM4[8139]<=16'd57285;
ROM1[8140]<=16'd4861; ROM2[8140]<=16'd0; ROM3[8140]<=16'd23755; ROM4[8140]<=16'd57271;
ROM1[8141]<=16'd4850; ROM2[8141]<=16'd0; ROM3[8141]<=16'd23753; ROM4[8141]<=16'd57272;
ROM1[8142]<=16'd4845; ROM2[8142]<=16'd0; ROM3[8142]<=16'd23769; ROM4[8142]<=16'd57288;
ROM1[8143]<=16'd4828; ROM2[8143]<=16'd0; ROM3[8143]<=16'd23782; ROM4[8143]<=16'd57291;
ROM1[8144]<=16'd4819; ROM2[8144]<=16'd0; ROM3[8144]<=16'd23794; ROM4[8144]<=16'd57298;
ROM1[8145]<=16'd4809; ROM2[8145]<=16'd0; ROM3[8145]<=16'd23798; ROM4[8145]<=16'd57299;
ROM1[8146]<=16'd4809; ROM2[8146]<=16'd0; ROM3[8146]<=16'd23793; ROM4[8146]<=16'd57297;
ROM1[8147]<=16'd4824; ROM2[8147]<=16'd0; ROM3[8147]<=16'd23774; ROM4[8147]<=16'd57289;
ROM1[8148]<=16'd4845; ROM2[8148]<=16'd0; ROM3[8148]<=16'd23755; ROM4[8148]<=16'd57280;
ROM1[8149]<=16'd4851; ROM2[8149]<=16'd0; ROM3[8149]<=16'd23754; ROM4[8149]<=16'd57281;
ROM1[8150]<=16'd4838; ROM2[8150]<=16'd0; ROM3[8150]<=16'd23760; ROM4[8150]<=16'd57286;
ROM1[8151]<=16'd4823; ROM2[8151]<=16'd0; ROM3[8151]<=16'd23772; ROM4[8151]<=16'd57287;
ROM1[8152]<=16'd4826; ROM2[8152]<=16'd0; ROM3[8152]<=16'd23794; ROM4[8152]<=16'd57300;
ROM1[8153]<=16'd4826; ROM2[8153]<=16'd0; ROM3[8153]<=16'd23812; ROM4[8153]<=16'd57313;
ROM1[8154]<=16'd4816; ROM2[8154]<=16'd0; ROM3[8154]<=16'd23800; ROM4[8154]<=16'd57299;
ROM1[8155]<=16'd4818; ROM2[8155]<=16'd0; ROM3[8155]<=16'd23772; ROM4[8155]<=16'd57278;
ROM1[8156]<=16'd4844; ROM2[8156]<=16'd0; ROM3[8156]<=16'd23751; ROM4[8156]<=16'd57268;
ROM1[8157]<=16'd4852; ROM2[8157]<=16'd0; ROM3[8157]<=16'd23734; ROM4[8157]<=16'd57262;
ROM1[8158]<=16'd4835; ROM2[8158]<=16'd0; ROM3[8158]<=16'd23734; ROM4[8158]<=16'd57261;
ROM1[8159]<=16'd4819; ROM2[8159]<=16'd0; ROM3[8159]<=16'd23750; ROM4[8159]<=16'd57264;
ROM1[8160]<=16'd4799; ROM2[8160]<=16'd0; ROM3[8160]<=16'd23747; ROM4[8160]<=16'd57260;
ROM1[8161]<=16'd4782; ROM2[8161]<=16'd0; ROM3[8161]<=16'd23754; ROM4[8161]<=16'd57257;
ROM1[8162]<=16'd4794; ROM2[8162]<=16'd0; ROM3[8162]<=16'd23773; ROM4[8162]<=16'd57273;
ROM1[8163]<=16'd4823; ROM2[8163]<=16'd0; ROM3[8163]<=16'd23779; ROM4[8163]<=16'd57287;
ROM1[8164]<=16'd4851; ROM2[8164]<=16'd0; ROM3[8164]<=16'd23766; ROM4[8164]<=16'd57282;
ROM1[8165]<=16'd4869; ROM2[8165]<=16'd0; ROM3[8165]<=16'd23752; ROM4[8165]<=16'd57275;
ROM1[8166]<=16'd4845; ROM2[8166]<=16'd0; ROM3[8166]<=16'd23734; ROM4[8166]<=16'd57255;
ROM1[8167]<=16'd4817; ROM2[8167]<=16'd0; ROM3[8167]<=16'd23726; ROM4[8167]<=16'd57239;
ROM1[8168]<=16'd4796; ROM2[8168]<=16'd0; ROM3[8168]<=16'd23733; ROM4[8168]<=16'd57234;
ROM1[8169]<=16'd4780; ROM2[8169]<=16'd0; ROM3[8169]<=16'd23733; ROM4[8169]<=16'd57229;
ROM1[8170]<=16'd4777; ROM2[8170]<=16'd0; ROM3[8170]<=16'd23738; ROM4[8170]<=16'd57228;
ROM1[8171]<=16'd4779; ROM2[8171]<=16'd0; ROM3[8171]<=16'd23731; ROM4[8171]<=16'd57227;
ROM1[8172]<=16'd4805; ROM2[8172]<=16'd0; ROM3[8172]<=16'd23717; ROM4[8172]<=16'd57227;
ROM1[8173]<=16'd4838; ROM2[8173]<=16'd0; ROM3[8173]<=16'd23712; ROM4[8173]<=16'd57235;
ROM1[8174]<=16'd4839; ROM2[8174]<=16'd0; ROM3[8174]<=16'd23717; ROM4[8174]<=16'd57239;
ROM1[8175]<=16'd4826; ROM2[8175]<=16'd0; ROM3[8175]<=16'd23721; ROM4[8175]<=16'd57242;
ROM1[8176]<=16'd4816; ROM2[8176]<=16'd0; ROM3[8176]<=16'd23733; ROM4[8176]<=16'd57249;
ROM1[8177]<=16'd4805; ROM2[8177]<=16'd0; ROM3[8177]<=16'd23745; ROM4[8177]<=16'd57255;
ROM1[8178]<=16'd4800; ROM2[8178]<=16'd0; ROM3[8178]<=16'd23758; ROM4[8178]<=16'd57268;
ROM1[8179]<=16'd4815; ROM2[8179]<=16'd0; ROM3[8179]<=16'd23781; ROM4[8179]<=16'd57283;
ROM1[8180]<=16'd4844; ROM2[8180]<=16'd0; ROM3[8180]<=16'd23787; ROM4[8180]<=16'd57293;
ROM1[8181]<=16'd4884; ROM2[8181]<=16'd0; ROM3[8181]<=16'd23778; ROM4[8181]<=16'd57301;
ROM1[8182]<=16'd4892; ROM2[8182]<=16'd0; ROM3[8182]<=16'd23775; ROM4[8182]<=16'd57299;
ROM1[8183]<=16'd4878; ROM2[8183]<=16'd0; ROM3[8183]<=16'd23783; ROM4[8183]<=16'd57302;
ROM1[8184]<=16'd4865; ROM2[8184]<=16'd0; ROM3[8184]<=16'd23799; ROM4[8184]<=16'd57313;
ROM1[8185]<=16'd4846; ROM2[8185]<=16'd0; ROM3[8185]<=16'd23801; ROM4[8185]<=16'd57302;
ROM1[8186]<=16'd4831; ROM2[8186]<=16'd0; ROM3[8186]<=16'd23808; ROM4[8186]<=16'd57305;
ROM1[8187]<=16'd4820; ROM2[8187]<=16'd0; ROM3[8187]<=16'd23807; ROM4[8187]<=16'd57302;
ROM1[8188]<=16'd4835; ROM2[8188]<=16'd0; ROM3[8188]<=16'd23801; ROM4[8188]<=16'd57298;
ROM1[8189]<=16'd4874; ROM2[8189]<=16'd0; ROM3[8189]<=16'd23799; ROM4[8189]<=16'd57310;
ROM1[8190]<=16'd4897; ROM2[8190]<=16'd0; ROM3[8190]<=16'd23790; ROM4[8190]<=16'd57304;
ROM1[8191]<=16'd4896; ROM2[8191]<=16'd0; ROM3[8191]<=16'd23790; ROM4[8191]<=16'd57303;
ROM1[8192]<=16'd4869; ROM2[8192]<=16'd0; ROM3[8192]<=16'd23790; ROM4[8192]<=16'd57300;
ROM1[8193]<=16'd4852; ROM2[8193]<=16'd0; ROM3[8193]<=16'd23803; ROM4[8193]<=16'd57305;
ROM1[8194]<=16'd4849; ROM2[8194]<=16'd0; ROM3[8194]<=16'd23814; ROM4[8194]<=16'd57316;
ROM1[8195]<=16'd4827; ROM2[8195]<=16'd0; ROM3[8195]<=16'd23804; ROM4[8195]<=16'd57300;
ROM1[8196]<=16'd4824; ROM2[8196]<=16'd0; ROM3[8196]<=16'd23789; ROM4[8196]<=16'd57285;
ROM1[8197]<=16'd4847; ROM2[8197]<=16'd0; ROM3[8197]<=16'd23771; ROM4[8197]<=16'd57279;
ROM1[8198]<=16'd4871; ROM2[8198]<=16'd0; ROM3[8198]<=16'd23753; ROM4[8198]<=16'd57272;
ROM1[8199]<=16'd4875; ROM2[8199]<=16'd0; ROM3[8199]<=16'd23758; ROM4[8199]<=16'd57277;
ROM1[8200]<=16'd4861; ROM2[8200]<=16'd0; ROM3[8200]<=16'd23767; ROM4[8200]<=16'd57276;
ROM1[8201]<=16'd4847; ROM2[8201]<=16'd0; ROM3[8201]<=16'd23782; ROM4[8201]<=16'd57282;
ROM1[8202]<=16'd4848; ROM2[8202]<=16'd0; ROM3[8202]<=16'd23807; ROM4[8202]<=16'd57300;
ROM1[8203]<=16'd4837; ROM2[8203]<=16'd0; ROM3[8203]<=16'd23811; ROM4[8203]<=16'd57304;
ROM1[8204]<=16'd4822; ROM2[8204]<=16'd0; ROM3[8204]<=16'd23800; ROM4[8204]<=16'd57294;
ROM1[8205]<=16'd4841; ROM2[8205]<=16'd0; ROM3[8205]<=16'd23796; ROM4[8205]<=16'd57294;
ROM1[8206]<=16'd4878; ROM2[8206]<=16'd0; ROM3[8206]<=16'd23785; ROM4[8206]<=16'd57295;
ROM1[8207]<=16'd4882; ROM2[8207]<=16'd0; ROM3[8207]<=16'd23768; ROM4[8207]<=16'd57292;
ROM1[8208]<=16'd4866; ROM2[8208]<=16'd0; ROM3[8208]<=16'd23771; ROM4[8208]<=16'd57295;
ROM1[8209]<=16'd4837; ROM2[8209]<=16'd0; ROM3[8209]<=16'd23769; ROM4[8209]<=16'd57286;
ROM1[8210]<=16'd4811; ROM2[8210]<=16'd0; ROM3[8210]<=16'd23765; ROM4[8210]<=16'd57275;
ROM1[8211]<=16'd4808; ROM2[8211]<=16'd0; ROM3[8211]<=16'd23784; ROM4[8211]<=16'd57283;
ROM1[8212]<=16'd4822; ROM2[8212]<=16'd0; ROM3[8212]<=16'd23795; ROM4[8212]<=16'd57297;
ROM1[8213]<=16'd4837; ROM2[8213]<=16'd0; ROM3[8213]<=16'd23784; ROM4[8213]<=16'd57293;
ROM1[8214]<=16'd4854; ROM2[8214]<=16'd0; ROM3[8214]<=16'd23764; ROM4[8214]<=16'd57282;
ROM1[8215]<=16'd4867; ROM2[8215]<=16'd0; ROM3[8215]<=16'd23755; ROM4[8215]<=16'd57276;
ROM1[8216]<=16'd4869; ROM2[8216]<=16'd0; ROM3[8216]<=16'd23772; ROM4[8216]<=16'd57289;
ROM1[8217]<=16'd4854; ROM2[8217]<=16'd0; ROM3[8217]<=16'd23788; ROM4[8217]<=16'd57297;
ROM1[8218]<=16'd4817; ROM2[8218]<=16'd0; ROM3[8218]<=16'd23774; ROM4[8218]<=16'd57279;
ROM1[8219]<=16'd4808; ROM2[8219]<=16'd0; ROM3[8219]<=16'd23779; ROM4[8219]<=16'd57282;
ROM1[8220]<=16'd4811; ROM2[8220]<=16'd0; ROM3[8220]<=16'd23789; ROM4[8220]<=16'd57293;
ROM1[8221]<=16'd4814; ROM2[8221]<=16'd0; ROM3[8221]<=16'd23786; ROM4[8221]<=16'd57290;
ROM1[8222]<=16'd4840; ROM2[8222]<=16'd0; ROM3[8222]<=16'd23784; ROM4[8222]<=16'd57289;
ROM1[8223]<=16'd4866; ROM2[8223]<=16'd0; ROM3[8223]<=16'd23769; ROM4[8223]<=16'd57287;
ROM1[8224]<=16'd4856; ROM2[8224]<=16'd0; ROM3[8224]<=16'd23760; ROM4[8224]<=16'd57277;
ROM1[8225]<=16'd4841; ROM2[8225]<=16'd0; ROM3[8225]<=16'd23764; ROM4[8225]<=16'd57275;
ROM1[8226]<=16'd4839; ROM2[8226]<=16'd0; ROM3[8226]<=16'd23780; ROM4[8226]<=16'd57290;
ROM1[8227]<=16'd4826; ROM2[8227]<=16'd0; ROM3[8227]<=16'd23786; ROM4[8227]<=16'd57292;
ROM1[8228]<=16'd4807; ROM2[8228]<=16'd0; ROM3[8228]<=16'd23788; ROM4[8228]<=16'd57289;
ROM1[8229]<=16'd4809; ROM2[8229]<=16'd0; ROM3[8229]<=16'd23789; ROM4[8229]<=16'd57287;
ROM1[8230]<=16'd4834; ROM2[8230]<=16'd0; ROM3[8230]<=16'd23783; ROM4[8230]<=16'd57286;
ROM1[8231]<=16'd4870; ROM2[8231]<=16'd0; ROM3[8231]<=16'd23771; ROM4[8231]<=16'd57289;
ROM1[8232]<=16'd4877; ROM2[8232]<=16'd0; ROM3[8232]<=16'd23764; ROM4[8232]<=16'd57287;
ROM1[8233]<=16'd4862; ROM2[8233]<=16'd0; ROM3[8233]<=16'd23766; ROM4[8233]<=16'd57284;
ROM1[8234]<=16'd4852; ROM2[8234]<=16'd0; ROM3[8234]<=16'd23778; ROM4[8234]<=16'd57294;
ROM1[8235]<=16'd4836; ROM2[8235]<=16'd0; ROM3[8235]<=16'd23784; ROM4[8235]<=16'd57291;
ROM1[8236]<=16'd4816; ROM2[8236]<=16'd0; ROM3[8236]<=16'd23778; ROM4[8236]<=16'd57278;
ROM1[8237]<=16'd4808; ROM2[8237]<=16'd0; ROM3[8237]<=16'd23772; ROM4[8237]<=16'd57270;
ROM1[8238]<=16'd4815; ROM2[8238]<=16'd0; ROM3[8238]<=16'd23766; ROM4[8238]<=16'd57263;
ROM1[8239]<=16'd4846; ROM2[8239]<=16'd0; ROM3[8239]<=16'd23754; ROM4[8239]<=16'd57264;
ROM1[8240]<=16'd4880; ROM2[8240]<=16'd0; ROM3[8240]<=16'd23758; ROM4[8240]<=16'd57274;
ROM1[8241]<=16'd4880; ROM2[8241]<=16'd0; ROM3[8241]<=16'd23769; ROM4[8241]<=16'd57280;
ROM1[8242]<=16'd4850; ROM2[8242]<=16'd0; ROM3[8242]<=16'd23764; ROM4[8242]<=16'd57270;
ROM1[8243]<=16'd4820; ROM2[8243]<=16'd0; ROM3[8243]<=16'd23762; ROM4[8243]<=16'd57259;
ROM1[8244]<=16'd4806; ROM2[8244]<=16'd0; ROM3[8244]<=16'd23772; ROM4[8244]<=16'd57263;
ROM1[8245]<=16'd4805; ROM2[8245]<=16'd0; ROM3[8245]<=16'd23793; ROM4[8245]<=16'd57280;
ROM1[8246]<=16'd4807; ROM2[8246]<=16'd0; ROM3[8246]<=16'd23795; ROM4[8246]<=16'd57282;
ROM1[8247]<=16'd4833; ROM2[8247]<=16'd0; ROM3[8247]<=16'd23786; ROM4[8247]<=16'd57278;
ROM1[8248]<=16'd4869; ROM2[8248]<=16'd0; ROM3[8248]<=16'd23783; ROM4[8248]<=16'd57284;
ROM1[8249]<=16'd4850; ROM2[8249]<=16'd0; ROM3[8249]<=16'd23762; ROM4[8249]<=16'd57268;
ROM1[8250]<=16'd4837; ROM2[8250]<=16'd0; ROM3[8250]<=16'd23769; ROM4[8250]<=16'd57270;
ROM1[8251]<=16'd4836; ROM2[8251]<=16'd0; ROM3[8251]<=16'd23797; ROM4[8251]<=16'd57290;
ROM1[8252]<=16'd4808; ROM2[8252]<=16'd0; ROM3[8252]<=16'd23788; ROM4[8252]<=16'd57282;
ROM1[8253]<=16'd4788; ROM2[8253]<=16'd0; ROM3[8253]<=16'd23782; ROM4[8253]<=16'd57272;
ROM1[8254]<=16'd4797; ROM2[8254]<=16'd0; ROM3[8254]<=16'd23786; ROM4[8254]<=16'd57280;
ROM1[8255]<=16'd4826; ROM2[8255]<=16'd0; ROM3[8255]<=16'd23783; ROM4[8255]<=16'd57289;
ROM1[8256]<=16'd4875; ROM2[8256]<=16'd0; ROM3[8256]<=16'd23784; ROM4[8256]<=16'd57303;
ROM1[8257]<=16'd4881; ROM2[8257]<=16'd0; ROM3[8257]<=16'd23773; ROM4[8257]<=16'd57299;
ROM1[8258]<=16'd4854; ROM2[8258]<=16'd0; ROM3[8258]<=16'd23760; ROM4[8258]<=16'd57283;
ROM1[8259]<=16'd4838; ROM2[8259]<=16'd0; ROM3[8259]<=16'd23767; ROM4[8259]<=16'd57285;
ROM1[8260]<=16'd4824; ROM2[8260]<=16'd0; ROM3[8260]<=16'd23772; ROM4[8260]<=16'd57287;
ROM1[8261]<=16'd4815; ROM2[8261]<=16'd0; ROM3[8261]<=16'd23785; ROM4[8261]<=16'd57291;
ROM1[8262]<=16'd4810; ROM2[8262]<=16'd0; ROM3[8262]<=16'd23786; ROM4[8262]<=16'd57288;
ROM1[8263]<=16'd4813; ROM2[8263]<=16'd0; ROM3[8263]<=16'd23771; ROM4[8263]<=16'd57278;
ROM1[8264]<=16'd4834; ROM2[8264]<=16'd0; ROM3[8264]<=16'd23753; ROM4[8264]<=16'd57266;
ROM1[8265]<=16'd4872; ROM2[8265]<=16'd0; ROM3[8265]<=16'd23756; ROM4[8265]<=16'd57283;
ROM1[8266]<=16'd4908; ROM2[8266]<=16'd0; ROM3[8266]<=16'd23802; ROM4[8266]<=16'd57331;
ROM1[8267]<=16'd4881; ROM2[8267]<=16'd0; ROM3[8267]<=16'd23805; ROM4[8267]<=16'd57324;
ROM1[8268]<=16'd4839; ROM2[8268]<=16'd0; ROM3[8268]<=16'd23786; ROM4[8268]<=16'd57297;
ROM1[8269]<=16'd4823; ROM2[8269]<=16'd0; ROM3[8269]<=16'd23792; ROM4[8269]<=16'd57300;
ROM1[8270]<=16'd4805; ROM2[8270]<=16'd0; ROM3[8270]<=16'd23788; ROM4[8270]<=16'd57293;
ROM1[8271]<=16'd4815; ROM2[8271]<=16'd0; ROM3[8271]<=16'd23786; ROM4[8271]<=16'd57295;
ROM1[8272]<=16'd4854; ROM2[8272]<=16'd0; ROM3[8272]<=16'd23789; ROM4[8272]<=16'd57309;
ROM1[8273]<=16'd4883; ROM2[8273]<=16'd0; ROM3[8273]<=16'd23783; ROM4[8273]<=16'd57312;
ROM1[8274]<=16'd4874; ROM2[8274]<=16'd0; ROM3[8274]<=16'd23774; ROM4[8274]<=16'd57304;
ROM1[8275]<=16'd4857; ROM2[8275]<=16'd0; ROM3[8275]<=16'd23775; ROM4[8275]<=16'd57300;
ROM1[8276]<=16'd4840; ROM2[8276]<=16'd0; ROM3[8276]<=16'd23784; ROM4[8276]<=16'd57300;
ROM1[8277]<=16'd4823; ROM2[8277]<=16'd0; ROM3[8277]<=16'd23785; ROM4[8277]<=16'd57297;
ROM1[8278]<=16'd4809; ROM2[8278]<=16'd0; ROM3[8278]<=16'd23787; ROM4[8278]<=16'd57298;
ROM1[8279]<=16'd4815; ROM2[8279]<=16'd0; ROM3[8279]<=16'd23791; ROM4[8279]<=16'd57303;
ROM1[8280]<=16'd4839; ROM2[8280]<=16'd0; ROM3[8280]<=16'd23785; ROM4[8280]<=16'd57304;
ROM1[8281]<=16'd4872; ROM2[8281]<=16'd0; ROM3[8281]<=16'd23770; ROM4[8281]<=16'd57300;
ROM1[8282]<=16'd4870; ROM2[8282]<=16'd0; ROM3[8282]<=16'd23752; ROM4[8282]<=16'd57288;
ROM1[8283]<=16'd4850; ROM2[8283]<=16'd0; ROM3[8283]<=16'd23749; ROM4[8283]<=16'd57279;
ROM1[8284]<=16'd4834; ROM2[8284]<=16'd0; ROM3[8284]<=16'd23756; ROM4[8284]<=16'd57277;
ROM1[8285]<=16'd4819; ROM2[8285]<=16'd0; ROM3[8285]<=16'd23760; ROM4[8285]<=16'd57279;
ROM1[8286]<=16'd4815; ROM2[8286]<=16'd0; ROM3[8286]<=16'd23772; ROM4[8286]<=16'd57287;
ROM1[8287]<=16'd4813; ROM2[8287]<=16'd0; ROM3[8287]<=16'd23780; ROM4[8287]<=16'd57291;
ROM1[8288]<=16'd4821; ROM2[8288]<=16'd0; ROM3[8288]<=16'd23774; ROM4[8288]<=16'd57295;
ROM1[8289]<=16'd4856; ROM2[8289]<=16'd0; ROM3[8289]<=16'd23766; ROM4[8289]<=16'd57296;
ROM1[8290]<=16'd4886; ROM2[8290]<=16'd0; ROM3[8290]<=16'd23770; ROM4[8290]<=16'd57300;
ROM1[8291]<=16'd4880; ROM2[8291]<=16'd0; ROM3[8291]<=16'd23777; ROM4[8291]<=16'd57305;
ROM1[8292]<=16'd4869; ROM2[8292]<=16'd0; ROM3[8292]<=16'd23790; ROM4[8292]<=16'd57312;
ROM1[8293]<=16'd4862; ROM2[8293]<=16'd0; ROM3[8293]<=16'd23804; ROM4[8293]<=16'd57320;
ROM1[8294]<=16'd4842; ROM2[8294]<=16'd0; ROM3[8294]<=16'd23806; ROM4[8294]<=16'd57312;
ROM1[8295]<=16'd4835; ROM2[8295]<=16'd0; ROM3[8295]<=16'd23812; ROM4[8295]<=16'd57312;
ROM1[8296]<=16'd4847; ROM2[8296]<=16'd0; ROM3[8296]<=16'd23812; ROM4[8296]<=16'd57312;
ROM1[8297]<=16'd4871; ROM2[8297]<=16'd0; ROM3[8297]<=16'd23808; ROM4[8297]<=16'd57310;
ROM1[8298]<=16'd4895; ROM2[8298]<=16'd0; ROM3[8298]<=16'd23795; ROM4[8298]<=16'd57313;
ROM1[8299]<=16'd4885; ROM2[8299]<=16'd0; ROM3[8299]<=16'd23781; ROM4[8299]<=16'd57304;
ROM1[8300]<=16'd4863; ROM2[8300]<=16'd0; ROM3[8300]<=16'd23779; ROM4[8300]<=16'd57296;
ROM1[8301]<=16'd4840; ROM2[8301]<=16'd0; ROM3[8301]<=16'd23777; ROM4[8301]<=16'd57293;
ROM1[8302]<=16'd4826; ROM2[8302]<=16'd0; ROM3[8302]<=16'd23778; ROM4[8302]<=16'd57291;
ROM1[8303]<=16'd4817; ROM2[8303]<=16'd0; ROM3[8303]<=16'd23786; ROM4[8303]<=16'd57296;
ROM1[8304]<=16'd4820; ROM2[8304]<=16'd0; ROM3[8304]<=16'd23791; ROM4[8304]<=16'd57304;
ROM1[8305]<=16'd4847; ROM2[8305]<=16'd0; ROM3[8305]<=16'd23792; ROM4[8305]<=16'd57312;
ROM1[8306]<=16'd4898; ROM2[8306]<=16'd0; ROM3[8306]<=16'd23802; ROM4[8306]<=16'd57334;
ROM1[8307]<=16'd4909; ROM2[8307]<=16'd0; ROM3[8307]<=16'd23793; ROM4[8307]<=16'd57333;
ROM1[8308]<=16'd4872; ROM2[8308]<=16'd0; ROM3[8308]<=16'd23771; ROM4[8308]<=16'd57306;
ROM1[8309]<=16'd4850; ROM2[8309]<=16'd0; ROM3[8309]<=16'd23776; ROM4[8309]<=16'd57302;
ROM1[8310]<=16'd4827; ROM2[8310]<=16'd0; ROM3[8310]<=16'd23779; ROM4[8310]<=16'd57296;
ROM1[8311]<=16'd4793; ROM2[8311]<=16'd0; ROM3[8311]<=16'd23769; ROM4[8311]<=16'd57278;
ROM1[8312]<=16'd4792; ROM2[8312]<=16'd0; ROM3[8312]<=16'd23773; ROM4[8312]<=16'd57283;
ROM1[8313]<=16'd4810; ROM2[8313]<=16'd0; ROM3[8313]<=16'd23770; ROM4[8313]<=16'd57284;
ROM1[8314]<=16'd4842; ROM2[8314]<=16'd0; ROM3[8314]<=16'd23756; ROM4[8314]<=16'd57277;
ROM1[8315]<=16'd4881; ROM2[8315]<=16'd0; ROM3[8315]<=16'd23761; ROM4[8315]<=16'd57293;
ROM1[8316]<=16'd4887; ROM2[8316]<=16'd0; ROM3[8316]<=16'd23780; ROM4[8316]<=16'd57310;
ROM1[8317]<=16'd4858; ROM2[8317]<=16'd0; ROM3[8317]<=16'd23781; ROM4[8317]<=16'd57304;
ROM1[8318]<=16'd4834; ROM2[8318]<=16'd0; ROM3[8318]<=16'd23776; ROM4[8318]<=16'd57292;
ROM1[8319]<=16'd4828; ROM2[8319]<=16'd0; ROM3[8319]<=16'd23786; ROM4[8319]<=16'd57296;
ROM1[8320]<=16'd4826; ROM2[8320]<=16'd0; ROM3[8320]<=16'd23786; ROM4[8320]<=16'd57300;
ROM1[8321]<=16'd4836; ROM2[8321]<=16'd0; ROM3[8321]<=16'd23779; ROM4[8321]<=16'd57295;
ROM1[8322]<=16'd4851; ROM2[8322]<=16'd0; ROM3[8322]<=16'd23761; ROM4[8322]<=16'd57285;
ROM1[8323]<=16'd4871; ROM2[8323]<=16'd0; ROM3[8323]<=16'd23747; ROM4[8323]<=16'd57281;
ROM1[8324]<=16'd4867; ROM2[8324]<=16'd0; ROM3[8324]<=16'd23745; ROM4[8324]<=16'd57279;
ROM1[8325]<=16'd4846; ROM2[8325]<=16'd0; ROM3[8325]<=16'd23748; ROM4[8325]<=16'd57277;
ROM1[8326]<=16'd4838; ROM2[8326]<=16'd0; ROM3[8326]<=16'd23760; ROM4[8326]<=16'd57284;
ROM1[8327]<=16'd4835; ROM2[8327]<=16'd0; ROM3[8327]<=16'd23774; ROM4[8327]<=16'd57288;
ROM1[8328]<=16'd4829; ROM2[8328]<=16'd0; ROM3[8328]<=16'd23789; ROM4[8328]<=16'd57294;
ROM1[8329]<=16'd4828; ROM2[8329]<=16'd0; ROM3[8329]<=16'd23788; ROM4[8329]<=16'd57296;
ROM1[8330]<=16'd4841; ROM2[8330]<=16'd0; ROM3[8330]<=16'd23774; ROM4[8330]<=16'd57290;
ROM1[8331]<=16'd4855; ROM2[8331]<=16'd0; ROM3[8331]<=16'd23745; ROM4[8331]<=16'd57274;
ROM1[8332]<=16'd4855; ROM2[8332]<=16'd0; ROM3[8332]<=16'd23725; ROM4[8332]<=16'd57260;
ROM1[8333]<=16'd4843; ROM2[8333]<=16'd0; ROM3[8333]<=16'd23727; ROM4[8333]<=16'd57259;
ROM1[8334]<=16'd4830; ROM2[8334]<=16'd0; ROM3[8334]<=16'd23743; ROM4[8334]<=16'd57268;
ROM1[8335]<=16'd4833; ROM2[8335]<=16'd0; ROM3[8335]<=16'd23764; ROM4[8335]<=16'd57285;
ROM1[8336]<=16'd4806; ROM2[8336]<=16'd0; ROM3[8336]<=16'd23768; ROM4[8336]<=16'd57280;
ROM1[8337]<=16'd4788; ROM2[8337]<=16'd0; ROM3[8337]<=16'd23754; ROM4[8337]<=16'd57264;
ROM1[8338]<=16'd4799; ROM2[8338]<=16'd0; ROM3[8338]<=16'd23740; ROM4[8338]<=16'd57258;
ROM1[8339]<=16'd4827; ROM2[8339]<=16'd0; ROM3[8339]<=16'd23733; ROM4[8339]<=16'd57261;
ROM1[8340]<=16'd4858; ROM2[8340]<=16'd0; ROM3[8340]<=16'd23734; ROM4[8340]<=16'd57271;
ROM1[8341]<=16'd4875; ROM2[8341]<=16'd0; ROM3[8341]<=16'd23767; ROM4[8341]<=16'd57299;
ROM1[8342]<=16'd4853; ROM2[8342]<=16'd0; ROM3[8342]<=16'd23779; ROM4[8342]<=16'd57302;
ROM1[8343]<=16'd4819; ROM2[8343]<=16'd0; ROM3[8343]<=16'd23764; ROM4[8343]<=16'd57282;
ROM1[8344]<=16'd4799; ROM2[8344]<=16'd0; ROM3[8344]<=16'd23765; ROM4[8344]<=16'd57275;
ROM1[8345]<=16'd4777; ROM2[8345]<=16'd0; ROM3[8345]<=16'd23760; ROM4[8345]<=16'd57264;
ROM1[8346]<=16'd4779; ROM2[8346]<=16'd0; ROM3[8346]<=16'd23753; ROM4[8346]<=16'd57259;
ROM1[8347]<=16'd4817; ROM2[8347]<=16'd0; ROM3[8347]<=16'd23754; ROM4[8347]<=16'd57269;
ROM1[8348]<=16'd4850; ROM2[8348]<=16'd0; ROM3[8348]<=16'd23744; ROM4[8348]<=16'd57272;
ROM1[8349]<=16'd4857; ROM2[8349]<=16'd0; ROM3[8349]<=16'd23746; ROM4[8349]<=16'd57278;
ROM1[8350]<=16'd4867; ROM2[8350]<=16'd0; ROM3[8350]<=16'd23778; ROM4[8350]<=16'd57303;
ROM1[8351]<=16'd4841; ROM2[8351]<=16'd0; ROM3[8351]<=16'd23779; ROM4[8351]<=16'd57298;
ROM1[8352]<=16'd4802; ROM2[8352]<=16'd0; ROM3[8352]<=16'd23761; ROM4[8352]<=16'd57276;
ROM1[8353]<=16'd4787; ROM2[8353]<=16'd0; ROM3[8353]<=16'd23758; ROM4[8353]<=16'd57268;
ROM1[8354]<=16'd4774; ROM2[8354]<=16'd0; ROM3[8354]<=16'd23737; ROM4[8354]<=16'd57251;
ROM1[8355]<=16'd4799; ROM2[8355]<=16'd0; ROM3[8355]<=16'd23733; ROM4[8355]<=16'd57253;
ROM1[8356]<=16'd4849; ROM2[8356]<=16'd0; ROM3[8356]<=16'd23743; ROM4[8356]<=16'd57272;
ROM1[8357]<=16'd4853; ROM2[8357]<=16'd0; ROM3[8357]<=16'd23737; ROM4[8357]<=16'd57270;
ROM1[8358]<=16'd4840; ROM2[8358]<=16'd0; ROM3[8358]<=16'd23743; ROM4[8358]<=16'd57265;
ROM1[8359]<=16'd4839; ROM2[8359]<=16'd0; ROM3[8359]<=16'd23768; ROM4[8359]<=16'd57281;
ROM1[8360]<=16'd4829; ROM2[8360]<=16'd0; ROM3[8360]<=16'd23773; ROM4[8360]<=16'd57282;
ROM1[8361]<=16'd4800; ROM2[8361]<=16'd0; ROM3[8361]<=16'd23762; ROM4[8361]<=16'd57266;
ROM1[8362]<=16'd4807; ROM2[8362]<=16'd0; ROM3[8362]<=16'd23776; ROM4[8362]<=16'd57281;
ROM1[8363]<=16'd4824; ROM2[8363]<=16'd0; ROM3[8363]<=16'd23773; ROM4[8363]<=16'd57283;
ROM1[8364]<=16'd4846; ROM2[8364]<=16'd0; ROM3[8364]<=16'd23758; ROM4[8364]<=16'd57274;
ROM1[8365]<=16'd4871; ROM2[8365]<=16'd0; ROM3[8365]<=16'd23751; ROM4[8365]<=16'd57279;
ROM1[8366]<=16'd4864; ROM2[8366]<=16'd0; ROM3[8366]<=16'd23754; ROM4[8366]<=16'd57277;
ROM1[8367]<=16'd4847; ROM2[8367]<=16'd0; ROM3[8367]<=16'd23763; ROM4[8367]<=16'd57277;
ROM1[8368]<=16'd4829; ROM2[8368]<=16'd0; ROM3[8368]<=16'd23766; ROM4[8368]<=16'd57278;
ROM1[8369]<=16'd4816; ROM2[8369]<=16'd0; ROM3[8369]<=16'd23773; ROM4[8369]<=16'd57275;
ROM1[8370]<=16'd4786; ROM2[8370]<=16'd0; ROM3[8370]<=16'd23752; ROM4[8370]<=16'd57255;
ROM1[8371]<=16'd4779; ROM2[8371]<=16'd0; ROM3[8371]<=16'd23736; ROM4[8371]<=16'd57243;
ROM1[8372]<=16'd4814; ROM2[8372]<=16'd0; ROM3[8372]<=16'd23733; ROM4[8372]<=16'd57245;
ROM1[8373]<=16'd4840; ROM2[8373]<=16'd0; ROM3[8373]<=16'd23724; ROM4[8373]<=16'd57245;
ROM1[8374]<=16'd4833; ROM2[8374]<=16'd0; ROM3[8374]<=16'd23723; ROM4[8374]<=16'd57244;
ROM1[8375]<=16'd4821; ROM2[8375]<=16'd0; ROM3[8375]<=16'd23735; ROM4[8375]<=16'd57250;
ROM1[8376]<=16'd4823; ROM2[8376]<=16'd0; ROM3[8376]<=16'd23760; ROM4[8376]<=16'd57272;
ROM1[8377]<=16'd4810; ROM2[8377]<=16'd0; ROM3[8377]<=16'd23763; ROM4[8377]<=16'd57272;
ROM1[8378]<=16'd4792; ROM2[8378]<=16'd0; ROM3[8378]<=16'd23763; ROM4[8378]<=16'd57268;
ROM1[8379]<=16'd4785; ROM2[8379]<=16'd0; ROM3[8379]<=16'd23756; ROM4[8379]<=16'd57261;
ROM1[8380]<=16'd4786; ROM2[8380]<=16'd0; ROM3[8380]<=16'd23731; ROM4[8380]<=16'd57242;
ROM1[8381]<=16'd4813; ROM2[8381]<=16'd0; ROM3[8381]<=16'd23716; ROM4[8381]<=16'd57241;
ROM1[8382]<=16'd4829; ROM2[8382]<=16'd0; ROM3[8382]<=16'd23720; ROM4[8382]<=16'd57250;
ROM1[8383]<=16'd4818; ROM2[8383]<=16'd0; ROM3[8383]<=16'd23723; ROM4[8383]<=16'd57249;
ROM1[8384]<=16'd4804; ROM2[8384]<=16'd0; ROM3[8384]<=16'd23732; ROM4[8384]<=16'd57255;
ROM1[8385]<=16'd4798; ROM2[8385]<=16'd0; ROM3[8385]<=16'd23746; ROM4[8385]<=16'd57260;
ROM1[8386]<=16'd4784; ROM2[8386]<=16'd0; ROM3[8386]<=16'd23748; ROM4[8386]<=16'd57256;
ROM1[8387]<=16'd4779; ROM2[8387]<=16'd0; ROM3[8387]<=16'd23747; ROM4[8387]<=16'd57254;
ROM1[8388]<=16'd4792; ROM2[8388]<=16'd0; ROM3[8388]<=16'd23746; ROM4[8388]<=16'd57254;
ROM1[8389]<=16'd4829; ROM2[8389]<=16'd0; ROM3[8389]<=16'd23738; ROM4[8389]<=16'd57259;
ROM1[8390]<=16'd4852; ROM2[8390]<=16'd0; ROM3[8390]<=16'd23728; ROM4[8390]<=16'd57257;
ROM1[8391]<=16'd4846; ROM2[8391]<=16'd0; ROM3[8391]<=16'd23734; ROM4[8391]<=16'd57258;
ROM1[8392]<=16'd4824; ROM2[8392]<=16'd0; ROM3[8392]<=16'd23735; ROM4[8392]<=16'd57253;
ROM1[8393]<=16'd4805; ROM2[8393]<=16'd0; ROM3[8393]<=16'd23743; ROM4[8393]<=16'd57253;
ROM1[8394]<=16'd4788; ROM2[8394]<=16'd0; ROM3[8394]<=16'd23749; ROM4[8394]<=16'd57252;
ROM1[8395]<=16'd4779; ROM2[8395]<=16'd0; ROM3[8395]<=16'd23756; ROM4[8395]<=16'd57251;
ROM1[8396]<=16'd4805; ROM2[8396]<=16'd0; ROM3[8396]<=16'd23778; ROM4[8396]<=16'd57274;
ROM1[8397]<=16'd4841; ROM2[8397]<=16'd0; ROM3[8397]<=16'd23781; ROM4[8397]<=16'd57286;
ROM1[8398]<=16'd4854; ROM2[8398]<=16'd0; ROM3[8398]<=16'd23756; ROM4[8398]<=16'd57275;
ROM1[8399]<=16'd4837; ROM2[8399]<=16'd0; ROM3[8399]<=16'd23740; ROM4[8399]<=16'd57264;
ROM1[8400]<=16'd4820; ROM2[8400]<=16'd0; ROM3[8400]<=16'd23747; ROM4[8400]<=16'd57262;
ROM1[8401]<=16'd4812; ROM2[8401]<=16'd0; ROM3[8401]<=16'd23761; ROM4[8401]<=16'd57269;
ROM1[8402]<=16'd4809; ROM2[8402]<=16'd0; ROM3[8402]<=16'd23776; ROM4[8402]<=16'd57283;
ROM1[8403]<=16'd4813; ROM2[8403]<=16'd0; ROM3[8403]<=16'd23800; ROM4[8403]<=16'd57301;
ROM1[8404]<=16'd4831; ROM2[8404]<=16'd0; ROM3[8404]<=16'd23810; ROM4[8404]<=16'd57316;
ROM1[8405]<=16'd4831; ROM2[8405]<=16'd0; ROM3[8405]<=16'd23780; ROM4[8405]<=16'd57294;
ROM1[8406]<=16'd4850; ROM2[8406]<=16'd0; ROM3[8406]<=16'd23753; ROM4[8406]<=16'd57276;
ROM1[8407]<=16'd4861; ROM2[8407]<=16'd0; ROM3[8407]<=16'd23747; ROM4[8407]<=16'd57274;
ROM1[8408]<=16'd4838; ROM2[8408]<=16'd0; ROM3[8408]<=16'd23745; ROM4[8408]<=16'd57268;
ROM1[8409]<=16'd4824; ROM2[8409]<=16'd0; ROM3[8409]<=16'd23763; ROM4[8409]<=16'd57279;
ROM1[8410]<=16'd4823; ROM2[8410]<=16'd0; ROM3[8410]<=16'd23783; ROM4[8410]<=16'd57294;
ROM1[8411]<=16'd4803; ROM2[8411]<=16'd0; ROM3[8411]<=16'd23785; ROM4[8411]<=16'd57288;
ROM1[8412]<=16'd4790; ROM2[8412]<=16'd0; ROM3[8412]<=16'd23773; ROM4[8412]<=16'd57276;
ROM1[8413]<=16'd4806; ROM2[8413]<=16'd0; ROM3[8413]<=16'd23763; ROM4[8413]<=16'd57269;
ROM1[8414]<=16'd4830; ROM2[8414]<=16'd0; ROM3[8414]<=16'd23750; ROM4[8414]<=16'd57266;
ROM1[8415]<=16'd4839; ROM2[8415]<=16'd0; ROM3[8415]<=16'd23731; ROM4[8415]<=16'd57263;
ROM1[8416]<=16'd4818; ROM2[8416]<=16'd0; ROM3[8416]<=16'd23725; ROM4[8416]<=16'd57252;
ROM1[8417]<=16'd4792; ROM2[8417]<=16'd0; ROM3[8417]<=16'd23730; ROM4[8417]<=16'd57248;
ROM1[8418]<=16'd4786; ROM2[8418]<=16'd0; ROM3[8418]<=16'd23738; ROM4[8418]<=16'd57254;
ROM1[8419]<=16'd4771; ROM2[8419]<=16'd0; ROM3[8419]<=16'd23741; ROM4[8419]<=16'd57251;
ROM1[8420]<=16'd4759; ROM2[8420]<=16'd0; ROM3[8420]<=16'd23737; ROM4[8420]<=16'd57245;
ROM1[8421]<=16'd4769; ROM2[8421]<=16'd0; ROM3[8421]<=16'd23732; ROM4[8421]<=16'd57243;
ROM1[8422]<=16'd4792; ROM2[8422]<=16'd0; ROM3[8422]<=16'd23724; ROM4[8422]<=16'd57242;
ROM1[8423]<=16'd4820; ROM2[8423]<=16'd0; ROM3[8423]<=16'd23712; ROM4[8423]<=16'd57239;
ROM1[8424]<=16'd4815; ROM2[8424]<=16'd0; ROM3[8424]<=16'd23711; ROM4[8424]<=16'd57236;
ROM1[8425]<=16'd4793; ROM2[8425]<=16'd0; ROM3[8425]<=16'd23712; ROM4[8425]<=16'd57233;
ROM1[8426]<=16'd4780; ROM2[8426]<=16'd0; ROM3[8426]<=16'd23715; ROM4[8426]<=16'd57233;
ROM1[8427]<=16'd4769; ROM2[8427]<=16'd0; ROM3[8427]<=16'd23716; ROM4[8427]<=16'd57230;
ROM1[8428]<=16'd4752; ROM2[8428]<=16'd0; ROM3[8428]<=16'd23716; ROM4[8428]<=16'd57225;
ROM1[8429]<=16'd4755; ROM2[8429]<=16'd0; ROM3[8429]<=16'd23717; ROM4[8429]<=16'd57224;
ROM1[8430]<=16'd4773; ROM2[8430]<=16'd0; ROM3[8430]<=16'd23712; ROM4[8430]<=16'd57227;
ROM1[8431]<=16'd4799; ROM2[8431]<=16'd0; ROM3[8431]<=16'd23697; ROM4[8431]<=16'd57226;
ROM1[8432]<=16'd4811; ROM2[8432]<=16'd0; ROM3[8432]<=16'd23694; ROM4[8432]<=16'd57228;
ROM1[8433]<=16'd4806; ROM2[8433]<=16'd0; ROM3[8433]<=16'd23709; ROM4[8433]<=16'd57241;
ROM1[8434]<=16'd4790; ROM2[8434]<=16'd0; ROM3[8434]<=16'd23716; ROM4[8434]<=16'd57236;
ROM1[8435]<=16'd4770; ROM2[8435]<=16'd0; ROM3[8435]<=16'd23720; ROM4[8435]<=16'd57229;
ROM1[8436]<=16'd4749; ROM2[8436]<=16'd0; ROM3[8436]<=16'd23722; ROM4[8436]<=16'd57227;
ROM1[8437]<=16'd4743; ROM2[8437]<=16'd0; ROM3[8437]<=16'd23719; ROM4[8437]<=16'd57226;
ROM1[8438]<=16'd4764; ROM2[8438]<=16'd0; ROM3[8438]<=16'd23722; ROM4[8438]<=16'd57235;
ROM1[8439]<=16'd4817; ROM2[8439]<=16'd0; ROM3[8439]<=16'd23734; ROM4[8439]<=16'd57258;
ROM1[8440]<=16'd4855; ROM2[8440]<=16'd0; ROM3[8440]<=16'd23750; ROM4[8440]<=16'd57282;
ROM1[8441]<=16'd4825; ROM2[8441]<=16'd0; ROM3[8441]<=16'd23735; ROM4[8441]<=16'd57265;
ROM1[8442]<=16'd4807; ROM2[8442]<=16'd0; ROM3[8442]<=16'd23749; ROM4[8442]<=16'd57267;
ROM1[8443]<=16'd4810; ROM2[8443]<=16'd0; ROM3[8443]<=16'd23775; ROM4[8443]<=16'd57286;
ROM1[8444]<=16'd4790; ROM2[8444]<=16'd0; ROM3[8444]<=16'd23761; ROM4[8444]<=16'd57273;
ROM1[8445]<=16'd4797; ROM2[8445]<=16'd0; ROM3[8445]<=16'd23767; ROM4[8445]<=16'd57278;
ROM1[8446]<=16'd4804; ROM2[8446]<=16'd0; ROM3[8446]<=16'd23755; ROM4[8446]<=16'd57269;
ROM1[8447]<=16'd4811; ROM2[8447]<=16'd0; ROM3[8447]<=16'd23730; ROM4[8447]<=16'd57248;
ROM1[8448]<=16'd4840; ROM2[8448]<=16'd0; ROM3[8448]<=16'd23725; ROM4[8448]<=16'd57253;
ROM1[8449]<=16'd4836; ROM2[8449]<=16'd0; ROM3[8449]<=16'd23727; ROM4[8449]<=16'd57253;
ROM1[8450]<=16'd4818; ROM2[8450]<=16'd0; ROM3[8450]<=16'd23734; ROM4[8450]<=16'd57252;
ROM1[8451]<=16'd4826; ROM2[8451]<=16'd0; ROM3[8451]<=16'd23753; ROM4[8451]<=16'd57269;
ROM1[8452]<=16'd4823; ROM2[8452]<=16'd0; ROM3[8452]<=16'd23766; ROM4[8452]<=16'd57277;
ROM1[8453]<=16'd4803; ROM2[8453]<=16'd0; ROM3[8453]<=16'd23769; ROM4[8453]<=16'd57267;
ROM1[8454]<=16'd4804; ROM2[8454]<=16'd0; ROM3[8454]<=16'd23766; ROM4[8454]<=16'd57266;
ROM1[8455]<=16'd4820; ROM2[8455]<=16'd0; ROM3[8455]<=16'd23751; ROM4[8455]<=16'd57264;
ROM1[8456]<=16'd4844; ROM2[8456]<=16'd0; ROM3[8456]<=16'd23734; ROM4[8456]<=16'd57254;
ROM1[8457]<=16'd4855; ROM2[8457]<=16'd0; ROM3[8457]<=16'd23731; ROM4[8457]<=16'd57253;
ROM1[8458]<=16'd4842; ROM2[8458]<=16'd0; ROM3[8458]<=16'd23737; ROM4[8458]<=16'd57259;
ROM1[8459]<=16'd4814; ROM2[8459]<=16'd0; ROM3[8459]<=16'd23742; ROM4[8459]<=16'd57252;
ROM1[8460]<=16'd4797; ROM2[8460]<=16'd0; ROM3[8460]<=16'd23749; ROM4[8460]<=16'd57254;
ROM1[8461]<=16'd4791; ROM2[8461]<=16'd0; ROM3[8461]<=16'd23761; ROM4[8461]<=16'd57266;
ROM1[8462]<=16'd4786; ROM2[8462]<=16'd0; ROM3[8462]<=16'd23765; ROM4[8462]<=16'd57269;
ROM1[8463]<=16'd4789; ROM2[8463]<=16'd0; ROM3[8463]<=16'd23752; ROM4[8463]<=16'd57263;
ROM1[8464]<=16'd4819; ROM2[8464]<=16'd0; ROM3[8464]<=16'd23740; ROM4[8464]<=16'd57263;
ROM1[8465]<=16'd4841; ROM2[8465]<=16'd0; ROM3[8465]<=16'd23733; ROM4[8465]<=16'd57270;
ROM1[8466]<=16'd4829; ROM2[8466]<=16'd0; ROM3[8466]<=16'd23731; ROM4[8466]<=16'd57273;
ROM1[8467]<=16'd4806; ROM2[8467]<=16'd0; ROM3[8467]<=16'd23731; ROM4[8467]<=16'd57268;
ROM1[8468]<=16'd4791; ROM2[8468]<=16'd0; ROM3[8468]<=16'd23732; ROM4[8468]<=16'd57266;
ROM1[8469]<=16'd4771; ROM2[8469]<=16'd0; ROM3[8469]<=16'd23732; ROM4[8469]<=16'd57259;
ROM1[8470]<=16'd4758; ROM2[8470]<=16'd0; ROM3[8470]<=16'd23734; ROM4[8470]<=16'd57256;
ROM1[8471]<=16'd4768; ROM2[8471]<=16'd0; ROM3[8471]<=16'd23730; ROM4[8471]<=16'd57255;
ROM1[8472]<=16'd4801; ROM2[8472]<=16'd0; ROM3[8472]<=16'd23724; ROM4[8472]<=16'd57261;
ROM1[8473]<=16'd4833; ROM2[8473]<=16'd0; ROM3[8473]<=16'd23718; ROM4[8473]<=16'd57267;
ROM1[8474]<=16'd4823; ROM2[8474]<=16'd0; ROM3[8474]<=16'd23708; ROM4[8474]<=16'd57255;
ROM1[8475]<=16'd4801; ROM2[8475]<=16'd0; ROM3[8475]<=16'd23705; ROM4[8475]<=16'd57245;
ROM1[8476]<=16'd4778; ROM2[8476]<=16'd0; ROM3[8476]<=16'd23707; ROM4[8476]<=16'd57234;
ROM1[8477]<=16'd4761; ROM2[8477]<=16'd0; ROM3[8477]<=16'd23707; ROM4[8477]<=16'd57225;
ROM1[8478]<=16'd4751; ROM2[8478]<=16'd0; ROM3[8478]<=16'd23712; ROM4[8478]<=16'd57226;
ROM1[8479]<=16'd4759; ROM2[8479]<=16'd0; ROM3[8479]<=16'd23722; ROM4[8479]<=16'd57232;
ROM1[8480]<=16'd4783; ROM2[8480]<=16'd0; ROM3[8480]<=16'd23721; ROM4[8480]<=16'd57234;
ROM1[8481]<=16'd4816; ROM2[8481]<=16'd0; ROM3[8481]<=16'd23707; ROM4[8481]<=16'd57236;
ROM1[8482]<=16'd4818; ROM2[8482]<=16'd0; ROM3[8482]<=16'd23703; ROM4[8482]<=16'd57230;
ROM1[8483]<=16'd4787; ROM2[8483]<=16'd0; ROM3[8483]<=16'd23696; ROM4[8483]<=16'd57215;
ROM1[8484]<=16'd4782; ROM2[8484]<=16'd0; ROM3[8484]<=16'd23716; ROM4[8484]<=16'd57229;
ROM1[8485]<=16'd4773; ROM2[8485]<=16'd0; ROM3[8485]<=16'd23729; ROM4[8485]<=16'd57235;
ROM1[8486]<=16'd4746; ROM2[8486]<=16'd0; ROM3[8486]<=16'd23718; ROM4[8486]<=16'd57217;
ROM1[8487]<=16'd4752; ROM2[8487]<=16'd0; ROM3[8487]<=16'd23722; ROM4[8487]<=16'd57222;
ROM1[8488]<=16'd4766; ROM2[8488]<=16'd0; ROM3[8488]<=16'd23716; ROM4[8488]<=16'd57222;
ROM1[8489]<=16'd4796; ROM2[8489]<=16'd0; ROM3[8489]<=16'd23705; ROM4[8489]<=16'd57221;
ROM1[8490]<=16'd4833; ROM2[8490]<=16'd0; ROM3[8490]<=16'd23713; ROM4[8490]<=16'd57241;
ROM1[8491]<=16'd4811; ROM2[8491]<=16'd0; ROM3[8491]<=16'd23704; ROM4[8491]<=16'd57236;
ROM1[8492]<=16'd4779; ROM2[8492]<=16'd0; ROM3[8492]<=16'd23699; ROM4[8492]<=16'd57225;
ROM1[8493]<=16'd4756; ROM2[8493]<=16'd0; ROM3[8493]<=16'd23698; ROM4[8493]<=16'd57218;
ROM1[8494]<=16'd4747; ROM2[8494]<=16'd0; ROM3[8494]<=16'd23707; ROM4[8494]<=16'd57224;
ROM1[8495]<=16'd4756; ROM2[8495]<=16'd0; ROM3[8495]<=16'd23721; ROM4[8495]<=16'd57236;
ROM1[8496]<=16'd4766; ROM2[8496]<=16'd0; ROM3[8496]<=16'd23719; ROM4[8496]<=16'd57236;
ROM1[8497]<=16'd4795; ROM2[8497]<=16'd0; ROM3[8497]<=16'd23714; ROM4[8497]<=16'd57238;
ROM1[8498]<=16'd4829; ROM2[8498]<=16'd0; ROM3[8498]<=16'd23705; ROM4[8498]<=16'd57238;
ROM1[8499]<=16'd4835; ROM2[8499]<=16'd0; ROM3[8499]<=16'd23709; ROM4[8499]<=16'd57249;
ROM1[8500]<=16'd4817; ROM2[8500]<=16'd0; ROM3[8500]<=16'd23716; ROM4[8500]<=16'd57252;
ROM1[8501]<=16'd4811; ROM2[8501]<=16'd0; ROM3[8501]<=16'd23732; ROM4[8501]<=16'd57258;
ROM1[8502]<=16'd4809; ROM2[8502]<=16'd0; ROM3[8502]<=16'd23750; ROM4[8502]<=16'd57270;
ROM1[8503]<=16'd4773; ROM2[8503]<=16'd0; ROM3[8503]<=16'd23735; ROM4[8503]<=16'd57249;
ROM1[8504]<=16'd4767; ROM2[8504]<=16'd0; ROM3[8504]<=16'd23722; ROM4[8504]<=16'd57235;
ROM1[8505]<=16'd4795; ROM2[8505]<=16'd0; ROM3[8505]<=16'd23716; ROM4[8505]<=16'd57239;
ROM1[8506]<=16'd4823; ROM2[8506]<=16'd0; ROM3[8506]<=16'd23705; ROM4[8506]<=16'd57235;
ROM1[8507]<=16'd4835; ROM2[8507]<=16'd0; ROM3[8507]<=16'd23708; ROM4[8507]<=16'd57239;
ROM1[8508]<=16'd4819; ROM2[8508]<=16'd0; ROM3[8508]<=16'd23712; ROM4[8508]<=16'd57240;
ROM1[8509]<=16'd4803; ROM2[8509]<=16'd0; ROM3[8509]<=16'd23724; ROM4[8509]<=16'd57246;
ROM1[8510]<=16'd4786; ROM2[8510]<=16'd0; ROM3[8510]<=16'd23731; ROM4[8510]<=16'd57245;
ROM1[8511]<=16'd4784; ROM2[8511]<=16'd0; ROM3[8511]<=16'd23751; ROM4[8511]<=16'd57256;
ROM1[8512]<=16'd4791; ROM2[8512]<=16'd0; ROM3[8512]<=16'd23762; ROM4[8512]<=16'd57267;
ROM1[8513]<=16'd4791; ROM2[8513]<=16'd0; ROM3[8513]<=16'd23739; ROM4[8513]<=16'd57253;
ROM1[8514]<=16'd4812; ROM2[8514]<=16'd0; ROM3[8514]<=16'd23716; ROM4[8514]<=16'd57243;
ROM1[8515]<=16'd4823; ROM2[8515]<=16'd0; ROM3[8515]<=16'd23699; ROM4[8515]<=16'd57232;
ROM1[8516]<=16'd4819; ROM2[8516]<=16'd0; ROM3[8516]<=16'd23702; ROM4[8516]<=16'd57230;
ROM1[8517]<=16'd4805; ROM2[8517]<=16'd0; ROM3[8517]<=16'd23711; ROM4[8517]<=16'd57229;
ROM1[8518]<=16'd4782; ROM2[8518]<=16'd0; ROM3[8518]<=16'd23711; ROM4[8518]<=16'd57225;
ROM1[8519]<=16'd4772; ROM2[8519]<=16'd0; ROM3[8519]<=16'd23719; ROM4[8519]<=16'd57227;
ROM1[8520]<=16'd4761; ROM2[8520]<=16'd0; ROM3[8520]<=16'd23720; ROM4[8520]<=16'd57226;
ROM1[8521]<=16'd4759; ROM2[8521]<=16'd0; ROM3[8521]<=16'd23705; ROM4[8521]<=16'd57215;
ROM1[8522]<=16'd4781; ROM2[8522]<=16'd0; ROM3[8522]<=16'd23686; ROM4[8522]<=16'd57205;
ROM1[8523]<=16'd4818; ROM2[8523]<=16'd0; ROM3[8523]<=16'd23685; ROM4[8523]<=16'd57217;
ROM1[8524]<=16'd4805; ROM2[8524]<=16'd0; ROM3[8524]<=16'd23682; ROM4[8524]<=16'd57212;
ROM1[8525]<=16'd4767; ROM2[8525]<=16'd0; ROM3[8525]<=16'd23673; ROM4[8525]<=16'd57198;
ROM1[8526]<=16'd4754; ROM2[8526]<=16'd0; ROM3[8526]<=16'd23686; ROM4[8526]<=16'd57203;
ROM1[8527]<=16'd4736; ROM2[8527]<=16'd0; ROM3[8527]<=16'd23686; ROM4[8527]<=16'd57199;
ROM1[8528]<=16'd4718; ROM2[8528]<=16'd0; ROM3[8528]<=16'd23683; ROM4[8528]<=16'd57194;
ROM1[8529]<=16'd4726; ROM2[8529]<=16'd0; ROM3[8529]<=16'd23689; ROM4[8529]<=16'd57198;
ROM1[8530]<=16'd4760; ROM2[8530]<=16'd0; ROM3[8530]<=16'd23695; ROM4[8530]<=16'd57211;
ROM1[8531]<=16'd4797; ROM2[8531]<=16'd0; ROM3[8531]<=16'd23692; ROM4[8531]<=16'd57222;
ROM1[8532]<=16'd4814; ROM2[8532]<=16'd0; ROM3[8532]<=16'd23700; ROM4[8532]<=16'd57234;
ROM1[8533]<=16'd4813; ROM2[8533]<=16'd0; ROM3[8533]<=16'd23723; ROM4[8533]<=16'd57249;
ROM1[8534]<=16'd4793; ROM2[8534]<=16'd0; ROM3[8534]<=16'd23732; ROM4[8534]<=16'd57251;
ROM1[8535]<=16'd4763; ROM2[8535]<=16'd0; ROM3[8535]<=16'd23721; ROM4[8535]<=16'd57228;
ROM1[8536]<=16'd4738; ROM2[8536]<=16'd0; ROM3[8536]<=16'd23713; ROM4[8536]<=16'd57214;
ROM1[8537]<=16'd4727; ROM2[8537]<=16'd0; ROM3[8537]<=16'd23702; ROM4[8537]<=16'd57204;
ROM1[8538]<=16'd4736; ROM2[8538]<=16'd0; ROM3[8538]<=16'd23688; ROM4[8538]<=16'd57196;
ROM1[8539]<=16'd4773; ROM2[8539]<=16'd0; ROM3[8539]<=16'd23681; ROM4[8539]<=16'd57202;
ROM1[8540]<=16'd4797; ROM2[8540]<=16'd0; ROM3[8540]<=16'd23677; ROM4[8540]<=16'd57209;
ROM1[8541]<=16'd4786; ROM2[8541]<=16'd0; ROM3[8541]<=16'd23677; ROM4[8541]<=16'd57212;
ROM1[8542]<=16'd4774; ROM2[8542]<=16'd0; ROM3[8542]<=16'd23687; ROM4[8542]<=16'd57214;
ROM1[8543]<=16'd4764; ROM2[8543]<=16'd0; ROM3[8543]<=16'd23701; ROM4[8543]<=16'd57221;
ROM1[8544]<=16'd4759; ROM2[8544]<=16'd0; ROM3[8544]<=16'd23723; ROM4[8544]<=16'd57236;
ROM1[8545]<=16'd4758; ROM2[8545]<=16'd0; ROM3[8545]<=16'd23734; ROM4[8545]<=16'd57241;
ROM1[8546]<=16'd4762; ROM2[8546]<=16'd0; ROM3[8546]<=16'd23720; ROM4[8546]<=16'd57233;
ROM1[8547]<=16'd4793; ROM2[8547]<=16'd0; ROM3[8547]<=16'd23711; ROM4[8547]<=16'd57239;
ROM1[8548]<=16'd4834; ROM2[8548]<=16'd0; ROM3[8548]<=16'd23714; ROM4[8548]<=16'd57254;
ROM1[8549]<=16'd4829; ROM2[8549]<=16'd0; ROM3[8549]<=16'd23714; ROM4[8549]<=16'd57257;
ROM1[8550]<=16'd4793; ROM2[8550]<=16'd0; ROM3[8550]<=16'd23700; ROM4[8550]<=16'd57240;
ROM1[8551]<=16'd4768; ROM2[8551]<=16'd0; ROM3[8551]<=16'd23697; ROM4[8551]<=16'd57224;
ROM1[8552]<=16'd4752; ROM2[8552]<=16'd0; ROM3[8552]<=16'd23693; ROM4[8552]<=16'd57218;
ROM1[8553]<=16'd4735; ROM2[8553]<=16'd0; ROM3[8553]<=16'd23695; ROM4[8553]<=16'd57214;
ROM1[8554]<=16'd4754; ROM2[8554]<=16'd0; ROM3[8554]<=16'd23710; ROM4[8554]<=16'd57225;
ROM1[8555]<=16'd4777; ROM2[8555]<=16'd0; ROM3[8555]<=16'd23698; ROM4[8555]<=16'd57224;
ROM1[8556]<=16'd4805; ROM2[8556]<=16'd0; ROM3[8556]<=16'd23679; ROM4[8556]<=16'd57218;
ROM1[8557]<=16'd4823; ROM2[8557]<=16'd0; ROM3[8557]<=16'd23680; ROM4[8557]<=16'd57226;
ROM1[8558]<=16'd4819; ROM2[8558]<=16'd0; ROM3[8558]<=16'd23698; ROM4[8558]<=16'd57239;
ROM1[8559]<=16'd4814; ROM2[8559]<=16'd0; ROM3[8559]<=16'd23727; ROM4[8559]<=16'd57260;
ROM1[8560]<=16'd4800; ROM2[8560]<=16'd0; ROM3[8560]<=16'd23736; ROM4[8560]<=16'd57263;
ROM1[8561]<=16'd4763; ROM2[8561]<=16'd0; ROM3[8561]<=16'd23722; ROM4[8561]<=16'd57237;
ROM1[8562]<=16'd4746; ROM2[8562]<=16'd0; ROM3[8562]<=16'd23707; ROM4[8562]<=16'd57224;
ROM1[8563]<=16'd4763; ROM2[8563]<=16'd0; ROM3[8563]<=16'd23697; ROM4[8563]<=16'd57226;
ROM1[8564]<=16'd4796; ROM2[8564]<=16'd0; ROM3[8564]<=16'd23684; ROM4[8564]<=16'd57223;
ROM1[8565]<=16'd4830; ROM2[8565]<=16'd0; ROM3[8565]<=16'd23690; ROM4[8565]<=16'd57240;
ROM1[8566]<=16'd4826; ROM2[8566]<=16'd0; ROM3[8566]<=16'd23702; ROM4[8566]<=16'd57249;
ROM1[8567]<=16'd4783; ROM2[8567]<=16'd0; ROM3[8567]<=16'd23686; ROM4[8567]<=16'd57226;
ROM1[8568]<=16'd4756; ROM2[8568]<=16'd0; ROM3[8568]<=16'd23681; ROM4[8568]<=16'd57213;
ROM1[8569]<=16'd4745; ROM2[8569]<=16'd0; ROM3[8569]<=16'd23691; ROM4[8569]<=16'd57216;
ROM1[8570]<=16'd4748; ROM2[8570]<=16'd0; ROM3[8570]<=16'd23704; ROM4[8570]<=16'd57226;
ROM1[8571]<=16'd4763; ROM2[8571]<=16'd0; ROM3[8571]<=16'd23709; ROM4[8571]<=16'd57230;
ROM1[8572]<=16'd4784; ROM2[8572]<=16'd0; ROM3[8572]<=16'd23696; ROM4[8572]<=16'd57222;
ROM1[8573]<=16'd4801; ROM2[8573]<=16'd0; ROM3[8573]<=16'd23678; ROM4[8573]<=16'd57215;
ROM1[8574]<=16'd4788; ROM2[8574]<=16'd0; ROM3[8574]<=16'd23676; ROM4[8574]<=16'd57208;
ROM1[8575]<=16'd4786; ROM2[8575]<=16'd0; ROM3[8575]<=16'd23709; ROM4[8575]<=16'd57230;
ROM1[8576]<=16'd4781; ROM2[8576]<=16'd0; ROM3[8576]<=16'd23728; ROM4[8576]<=16'd57245;
ROM1[8577]<=16'd4760; ROM2[8577]<=16'd0; ROM3[8577]<=16'd23717; ROM4[8577]<=16'd57231;
ROM1[8578]<=16'd4738; ROM2[8578]<=16'd0; ROM3[8578]<=16'd23713; ROM4[8578]<=16'd57224;
ROM1[8579]<=16'd4734; ROM2[8579]<=16'd0; ROM3[8579]<=16'd23704; ROM4[8579]<=16'd57219;
ROM1[8580]<=16'd4747; ROM2[8580]<=16'd0; ROM3[8580]<=16'd23687; ROM4[8580]<=16'd57209;
ROM1[8581]<=16'd4782; ROM2[8581]<=16'd0; ROM3[8581]<=16'd23683; ROM4[8581]<=16'd57218;
ROM1[8582]<=16'd4797; ROM2[8582]<=16'd0; ROM3[8582]<=16'd23687; ROM4[8582]<=16'd57224;
ROM1[8583]<=16'd4779; ROM2[8583]<=16'd0; ROM3[8583]<=16'd23688; ROM4[8583]<=16'd57218;
ROM1[8584]<=16'd4759; ROM2[8584]<=16'd0; ROM3[8584]<=16'd23693; ROM4[8584]<=16'd57216;
ROM1[8585]<=16'd4748; ROM2[8585]<=16'd0; ROM3[8585]<=16'd23696; ROM4[8585]<=16'd57215;
ROM1[8586]<=16'd4736; ROM2[8586]<=16'd0; ROM3[8586]<=16'd23697; ROM4[8586]<=16'd57215;
ROM1[8587]<=16'd4733; ROM2[8587]<=16'd0; ROM3[8587]<=16'd23698; ROM4[8587]<=16'd57216;
ROM1[8588]<=16'd4757; ROM2[8588]<=16'd0; ROM3[8588]<=16'd23701; ROM4[8588]<=16'd57222;
ROM1[8589]<=16'd4805; ROM2[8589]<=16'd0; ROM3[8589]<=16'd23710; ROM4[8589]<=16'd57236;
ROM1[8590]<=16'd4833; ROM2[8590]<=16'd0; ROM3[8590]<=16'd23721; ROM4[8590]<=16'd57249;
ROM1[8591]<=16'd4808; ROM2[8591]<=16'd0; ROM3[8591]<=16'd23709; ROM4[8591]<=16'd57231;
ROM1[8592]<=16'd4785; ROM2[8592]<=16'd0; ROM3[8592]<=16'd23712; ROM4[8592]<=16'd57229;
ROM1[8593]<=16'd4771; ROM2[8593]<=16'd0; ROM3[8593]<=16'd23722; ROM4[8593]<=16'd57236;
ROM1[8594]<=16'd4749; ROM2[8594]<=16'd0; ROM3[8594]<=16'd23718; ROM4[8594]<=16'd57227;
ROM1[8595]<=16'd4741; ROM2[8595]<=16'd0; ROM3[8595]<=16'd23718; ROM4[8595]<=16'd57226;
ROM1[8596]<=16'd4753; ROM2[8596]<=16'd0; ROM3[8596]<=16'd23720; ROM4[8596]<=16'd57229;
ROM1[8597]<=16'd4788; ROM2[8597]<=16'd0; ROM3[8597]<=16'd23719; ROM4[8597]<=16'd57236;
ROM1[8598]<=16'd4809; ROM2[8598]<=16'd0; ROM3[8598]<=16'd23694; ROM4[8598]<=16'd57225;
ROM1[8599]<=16'd4799; ROM2[8599]<=16'd0; ROM3[8599]<=16'd23683; ROM4[8599]<=16'd57215;
ROM1[8600]<=16'd4785; ROM2[8600]<=16'd0; ROM3[8600]<=16'd23686; ROM4[8600]<=16'd57216;
ROM1[8601]<=16'd4772; ROM2[8601]<=16'd0; ROM3[8601]<=16'd23691; ROM4[8601]<=16'd57216;
ROM1[8602]<=16'd4774; ROM2[8602]<=16'd0; ROM3[8602]<=16'd23705; ROM4[8602]<=16'd57232;
ROM1[8603]<=16'd4776; ROM2[8603]<=16'd0; ROM3[8603]<=16'd23717; ROM4[8603]<=16'd57243;
ROM1[8604]<=16'd4776; ROM2[8604]<=16'd0; ROM3[8604]<=16'd23714; ROM4[8604]<=16'd57238;
ROM1[8605]<=16'd4793; ROM2[8605]<=16'd0; ROM3[8605]<=16'd23701; ROM4[8605]<=16'd57234;
ROM1[8606]<=16'd4830; ROM2[8606]<=16'd0; ROM3[8606]<=16'd23693; ROM4[8606]<=16'd57239;
ROM1[8607]<=16'd4858; ROM2[8607]<=16'd0; ROM3[8607]<=16'd23710; ROM4[8607]<=16'd57260;
ROM1[8608]<=16'd4856; ROM2[8608]<=16'd0; ROM3[8608]<=16'd23726; ROM4[8608]<=16'd57273;
ROM1[8609]<=16'd4817; ROM2[8609]<=16'd0; ROM3[8609]<=16'd23720; ROM4[8609]<=16'd57257;
ROM1[8610]<=16'd4803; ROM2[8610]<=16'd0; ROM3[8610]<=16'd23727; ROM4[8610]<=16'd57260;
ROM1[8611]<=16'd4797; ROM2[8611]<=16'd0; ROM3[8611]<=16'd23736; ROM4[8611]<=16'd57266;
ROM1[8612]<=16'd4779; ROM2[8612]<=16'd0; ROM3[8612]<=16'd23718; ROM4[8612]<=16'd57252;
ROM1[8613]<=16'd4790; ROM2[8613]<=16'd0; ROM3[8613]<=16'd23697; ROM4[8613]<=16'd57246;
ROM1[8614]<=16'd4819; ROM2[8614]<=16'd0; ROM3[8614]<=16'd23683; ROM4[8614]<=16'd57238;
ROM1[8615]<=16'd4837; ROM2[8615]<=16'd0; ROM3[8615]<=16'd23677; ROM4[8615]<=16'd57241;
ROM1[8616]<=16'd4827; ROM2[8616]<=16'd0; ROM3[8616]<=16'd23678; ROM4[8616]<=16'd57243;
ROM1[8617]<=16'd4807; ROM2[8617]<=16'd0; ROM3[8617]<=16'd23683; ROM4[8617]<=16'd57239;
ROM1[8618]<=16'd4789; ROM2[8618]<=16'd0; ROM3[8618]<=16'd23688; ROM4[8618]<=16'd57237;
ROM1[8619]<=16'd4761; ROM2[8619]<=16'd0; ROM3[8619]<=16'd23680; ROM4[8619]<=16'd57222;
ROM1[8620]<=16'd4748; ROM2[8620]<=16'd0; ROM3[8620]<=16'd23682; ROM4[8620]<=16'd57217;
ROM1[8621]<=16'd4774; ROM2[8621]<=16'd0; ROM3[8621]<=16'd23698; ROM4[8621]<=16'd57229;
ROM1[8622]<=16'd4801; ROM2[8622]<=16'd0; ROM3[8622]<=16'd23693; ROM4[8622]<=16'd57229;
ROM1[8623]<=16'd4808; ROM2[8623]<=16'd0; ROM3[8623]<=16'd23669; ROM4[8623]<=16'd57217;
ROM1[8624]<=16'd4807; ROM2[8624]<=16'd0; ROM3[8624]<=16'd23674; ROM4[8624]<=16'd57220;
ROM1[8625]<=16'd4796; ROM2[8625]<=16'd0; ROM3[8625]<=16'd23690; ROM4[8625]<=16'd57226;
ROM1[8626]<=16'd4775; ROM2[8626]<=16'd0; ROM3[8626]<=16'd23700; ROM4[8626]<=16'd57230;
ROM1[8627]<=16'd4785; ROM2[8627]<=16'd0; ROM3[8627]<=16'd23731; ROM4[8627]<=16'd57257;
ROM1[8628]<=16'd4808; ROM2[8628]<=16'd0; ROM3[8628]<=16'd23766; ROM4[8628]<=16'd57288;
ROM1[8629]<=16'd4791; ROM2[8629]<=16'd0; ROM3[8629]<=16'd23744; ROM4[8629]<=16'd57270;
ROM1[8630]<=16'd4779; ROM2[8630]<=16'd0; ROM3[8630]<=16'd23702; ROM4[8630]<=16'd57231;
ROM1[8631]<=16'd4794; ROM2[8631]<=16'd0; ROM3[8631]<=16'd23673; ROM4[8631]<=16'd57213;
ROM1[8632]<=16'd4790; ROM2[8632]<=16'd0; ROM3[8632]<=16'd23657; ROM4[8632]<=16'd57199;
ROM1[8633]<=16'd4783; ROM2[8633]<=16'd0; ROM3[8633]<=16'd23667; ROM4[8633]<=16'd57203;
ROM1[8634]<=16'd4780; ROM2[8634]<=16'd0; ROM3[8634]<=16'd23691; ROM4[8634]<=16'd57224;
ROM1[8635]<=16'd4768; ROM2[8635]<=16'd0; ROM3[8635]<=16'd23698; ROM4[8635]<=16'd57220;
ROM1[8636]<=16'd4736; ROM2[8636]<=16'd0; ROM3[8636]<=16'd23691; ROM4[8636]<=16'd57207;
ROM1[8637]<=16'd4731; ROM2[8637]<=16'd0; ROM3[8637]<=16'd23701; ROM4[8637]<=16'd57212;
ROM1[8638]<=16'd4761; ROM2[8638]<=16'd0; ROM3[8638]<=16'd23709; ROM4[8638]<=16'd57222;
ROM1[8639]<=16'd4794; ROM2[8639]<=16'd0; ROM3[8639]<=16'd23703; ROM4[8639]<=16'd57222;
ROM1[8640]<=16'd4809; ROM2[8640]<=16'd0; ROM3[8640]<=16'd23700; ROM4[8640]<=16'd57222;
ROM1[8641]<=16'd4805; ROM2[8641]<=16'd0; ROM3[8641]<=16'd23708; ROM4[8641]<=16'd57229;
ROM1[8642]<=16'd4785; ROM2[8642]<=16'd0; ROM3[8642]<=16'd23715; ROM4[8642]<=16'd57230;
ROM1[8643]<=16'd4779; ROM2[8643]<=16'd0; ROM3[8643]<=16'd23733; ROM4[8643]<=16'd57238;
ROM1[8644]<=16'd4773; ROM2[8644]<=16'd0; ROM3[8644]<=16'd23742; ROM4[8644]<=16'd57240;
ROM1[8645]<=16'd4765; ROM2[8645]<=16'd0; ROM3[8645]<=16'd23741; ROM4[8645]<=16'd57237;
ROM1[8646]<=16'd4788; ROM2[8646]<=16'd0; ROM3[8646]<=16'd23744; ROM4[8646]<=16'd57250;
ROM1[8647]<=16'd4807; ROM2[8647]<=16'd0; ROM3[8647]<=16'd23724; ROM4[8647]<=16'd57243;
ROM1[8648]<=16'd4822; ROM2[8648]<=16'd0; ROM3[8648]<=16'd23702; ROM4[8648]<=16'd57229;
ROM1[8649]<=16'd4818; ROM2[8649]<=16'd0; ROM3[8649]<=16'd23696; ROM4[8649]<=16'd57227;
ROM1[8650]<=16'd4806; ROM2[8650]<=16'd0; ROM3[8650]<=16'd23705; ROM4[8650]<=16'd57231;
ROM1[8651]<=16'd4808; ROM2[8651]<=16'd0; ROM3[8651]<=16'd23729; ROM4[8651]<=16'd57250;
ROM1[8652]<=16'd4791; ROM2[8652]<=16'd0; ROM3[8652]<=16'd23730; ROM4[8652]<=16'd57248;
ROM1[8653]<=16'd4771; ROM2[8653]<=16'd0; ROM3[8653]<=16'd23726; ROM4[8653]<=16'd57241;
ROM1[8654]<=16'd4768; ROM2[8654]<=16'd0; ROM3[8654]<=16'd23721; ROM4[8654]<=16'd57236;
ROM1[8655]<=16'd4777; ROM2[8655]<=16'd0; ROM3[8655]<=16'd23694; ROM4[8655]<=16'd57217;
ROM1[8656]<=16'd4808; ROM2[8656]<=16'd0; ROM3[8656]<=16'd23680; ROM4[8656]<=16'd57219;
ROM1[8657]<=16'd4818; ROM2[8657]<=16'd0; ROM3[8657]<=16'd23684; ROM4[8657]<=16'd57225;
ROM1[8658]<=16'd4796; ROM2[8658]<=16'd0; ROM3[8658]<=16'd23680; ROM4[8658]<=16'd57216;
ROM1[8659]<=16'd4766; ROM2[8659]<=16'd0; ROM3[8659]<=16'd23680; ROM4[8659]<=16'd57210;
ROM1[8660]<=16'd4760; ROM2[8660]<=16'd0; ROM3[8660]<=16'd23694; ROM4[8660]<=16'd57219;
ROM1[8661]<=16'd4757; ROM2[8661]<=16'd0; ROM3[8661]<=16'd23712; ROM4[8661]<=16'd57230;
ROM1[8662]<=16'd4754; ROM2[8662]<=16'd0; ROM3[8662]<=16'd23717; ROM4[8662]<=16'd57232;
ROM1[8663]<=16'd4792; ROM2[8663]<=16'd0; ROM3[8663]<=16'd23736; ROM4[8663]<=16'd57258;
ROM1[8664]<=16'd4844; ROM2[8664]<=16'd0; ROM3[8664]<=16'd23748; ROM4[8664]<=16'd57283;
ROM1[8665]<=16'd4847; ROM2[8665]<=16'd0; ROM3[8665]<=16'd23723; ROM4[8665]<=16'd57269;
ROM1[8666]<=16'd4811; ROM2[8666]<=16'd0; ROM3[8666]<=16'd23700; ROM4[8666]<=16'd57242;
ROM1[8667]<=16'd4780; ROM2[8667]<=16'd0; ROM3[8667]<=16'd23694; ROM4[8667]<=16'd57227;
ROM1[8668]<=16'd4759; ROM2[8668]<=16'd0; ROM3[8668]<=16'd23696; ROM4[8668]<=16'd57220;
ROM1[8669]<=16'd4748; ROM2[8669]<=16'd0; ROM3[8669]<=16'd23709; ROM4[8669]<=16'd57224;
ROM1[8670]<=16'd4747; ROM2[8670]<=16'd0; ROM3[8670]<=16'd23722; ROM4[8670]<=16'd57236;
ROM1[8671]<=16'd4755; ROM2[8671]<=16'd0; ROM3[8671]<=16'd23719; ROM4[8671]<=16'd57237;
ROM1[8672]<=16'd4783; ROM2[8672]<=16'd0; ROM3[8672]<=16'd23705; ROM4[8672]<=16'd57232;
ROM1[8673]<=16'd4818; ROM2[8673]<=16'd0; ROM3[8673]<=16'd23700; ROM4[8673]<=16'd57240;
ROM1[8674]<=16'd4829; ROM2[8674]<=16'd0; ROM3[8674]<=16'd23712; ROM4[8674]<=16'd57256;
ROM1[8675]<=16'd4813; ROM2[8675]<=16'd0; ROM3[8675]<=16'd23719; ROM4[8675]<=16'd57258;
ROM1[8676]<=16'd4786; ROM2[8676]<=16'd0; ROM3[8676]<=16'd23715; ROM4[8676]<=16'd57250;
ROM1[8677]<=16'd4772; ROM2[8677]<=16'd0; ROM3[8677]<=16'd23718; ROM4[8677]<=16'd57250;
ROM1[8678]<=16'd4766; ROM2[8678]<=16'd0; ROM3[8678]<=16'd23728; ROM4[8678]<=16'd57257;
ROM1[8679]<=16'd4767; ROM2[8679]<=16'd0; ROM3[8679]<=16'd23724; ROM4[8679]<=16'd57257;
ROM1[8680]<=16'd4785; ROM2[8680]<=16'd0; ROM3[8680]<=16'd23710; ROM4[8680]<=16'd57253;
ROM1[8681]<=16'd4820; ROM2[8681]<=16'd0; ROM3[8681]<=16'd23698; ROM4[8681]<=16'd57253;
ROM1[8682]<=16'd4833; ROM2[8682]<=16'd0; ROM3[8682]<=16'd23696; ROM4[8682]<=16'd57251;
ROM1[8683]<=16'd4820; ROM2[8683]<=16'd0; ROM3[8683]<=16'd23701; ROM4[8683]<=16'd57253;
ROM1[8684]<=16'd4806; ROM2[8684]<=16'd0; ROM3[8684]<=16'd23711; ROM4[8684]<=16'd57256;
ROM1[8685]<=16'd4798; ROM2[8685]<=16'd0; ROM3[8685]<=16'd23723; ROM4[8685]<=16'd57261;
ROM1[8686]<=16'd4795; ROM2[8686]<=16'd0; ROM3[8686]<=16'd23741; ROM4[8686]<=16'd57274;
ROM1[8687]<=16'd4800; ROM2[8687]<=16'd0; ROM3[8687]<=16'd23753; ROM4[8687]<=16'd57282;
ROM1[8688]<=16'd4805; ROM2[8688]<=16'd0; ROM3[8688]<=16'd23739; ROM4[8688]<=16'd57273;
ROM1[8689]<=16'd4832; ROM2[8689]<=16'd0; ROM3[8689]<=16'd23726; ROM4[8689]<=16'd57266;
ROM1[8690]<=16'd4848; ROM2[8690]<=16'd0; ROM3[8690]<=16'd23716; ROM4[8690]<=16'd57263;
ROM1[8691]<=16'd4816; ROM2[8691]<=16'd0; ROM3[8691]<=16'd23695; ROM4[8691]<=16'd57240;
ROM1[8692]<=16'd4796; ROM2[8692]<=16'd0; ROM3[8692]<=16'd23699; ROM4[8692]<=16'd57237;
ROM1[8693]<=16'd4787; ROM2[8693]<=16'd0; ROM3[8693]<=16'd23710; ROM4[8693]<=16'd57242;
ROM1[8694]<=16'd4766; ROM2[8694]<=16'd0; ROM3[8694]<=16'd23713; ROM4[8694]<=16'd57239;
ROM1[8695]<=16'd4764; ROM2[8695]<=16'd0; ROM3[8695]<=16'd23720; ROM4[8695]<=16'd57240;
ROM1[8696]<=16'd4782; ROM2[8696]<=16'd0; ROM3[8696]<=16'd23727; ROM4[8696]<=16'd57248;
ROM1[8697]<=16'd4817; ROM2[8697]<=16'd0; ROM3[8697]<=16'd23729; ROM4[8697]<=16'd57257;
ROM1[8698]<=16'd4854; ROM2[8698]<=16'd0; ROM3[8698]<=16'd23730; ROM4[8698]<=16'd57265;
ROM1[8699]<=16'd4866; ROM2[8699]<=16'd0; ROM3[8699]<=16'd23744; ROM4[8699]<=16'd57283;
ROM1[8700]<=16'd4849; ROM2[8700]<=16'd0; ROM3[8700]<=16'd23753; ROM4[8700]<=16'd57285;
ROM1[8701]<=16'd4801; ROM2[8701]<=16'd0; ROM3[8701]<=16'd23734; ROM4[8701]<=16'd57258;
ROM1[8702]<=16'd4764; ROM2[8702]<=16'd0; ROM3[8702]<=16'd23716; ROM4[8702]<=16'd57235;
ROM1[8703]<=16'd4752; ROM2[8703]<=16'd0; ROM3[8703]<=16'd23719; ROM4[8703]<=16'd57233;
ROM1[8704]<=16'd4757; ROM2[8704]<=16'd0; ROM3[8704]<=16'd23717; ROM4[8704]<=16'd57233;
ROM1[8705]<=16'd4787; ROM2[8705]<=16'd0; ROM3[8705]<=16'd23710; ROM4[8705]<=16'd57240;
ROM1[8706]<=16'd4823; ROM2[8706]<=16'd0; ROM3[8706]<=16'd23701; ROM4[8706]<=16'd57244;
ROM1[8707]<=16'd4828; ROM2[8707]<=16'd0; ROM3[8707]<=16'd23702; ROM4[8707]<=16'd57247;
ROM1[8708]<=16'd4823; ROM2[8708]<=16'd0; ROM3[8708]<=16'd23716; ROM4[8708]<=16'd57252;
ROM1[8709]<=16'd4796; ROM2[8709]<=16'd0; ROM3[8709]<=16'd23717; ROM4[8709]<=16'd57242;
ROM1[8710]<=16'd4769; ROM2[8710]<=16'd0; ROM3[8710]<=16'd23707; ROM4[8710]<=16'd57231;
ROM1[8711]<=16'd4752; ROM2[8711]<=16'd0; ROM3[8711]<=16'd23706; ROM4[8711]<=16'd57225;
ROM1[8712]<=16'd4747; ROM2[8712]<=16'd0; ROM3[8712]<=16'd23708; ROM4[8712]<=16'd57227;
ROM1[8713]<=16'd4773; ROM2[8713]<=16'd0; ROM3[8713]<=16'd23708; ROM4[8713]<=16'd57239;
ROM1[8714]<=16'd4810; ROM2[8714]<=16'd0; ROM3[8714]<=16'd23702; ROM4[8714]<=16'd57242;
ROM1[8715]<=16'd4819; ROM2[8715]<=16'd0; ROM3[8715]<=16'd23685; ROM4[8715]<=16'd57233;
ROM1[8716]<=16'd4796; ROM2[8716]<=16'd0; ROM3[8716]<=16'd23668; ROM4[8716]<=16'd57220;
ROM1[8717]<=16'd4778; ROM2[8717]<=16'd0; ROM3[8717]<=16'd23671; ROM4[8717]<=16'd57220;
ROM1[8718]<=16'd4768; ROM2[8718]<=16'd0; ROM3[8718]<=16'd23682; ROM4[8718]<=16'd57226;
ROM1[8719]<=16'd4762; ROM2[8719]<=16'd0; ROM3[8719]<=16'd23692; ROM4[8719]<=16'd57234;
ROM1[8720]<=16'd4758; ROM2[8720]<=16'd0; ROM3[8720]<=16'd23701; ROM4[8720]<=16'd57238;
ROM1[8721]<=16'd4763; ROM2[8721]<=16'd0; ROM3[8721]<=16'd23697; ROM4[8721]<=16'd57236;
ROM1[8722]<=16'd4799; ROM2[8722]<=16'd0; ROM3[8722]<=16'd23692; ROM4[8722]<=16'd57240;
ROM1[8723]<=16'd4828; ROM2[8723]<=16'd0; ROM3[8723]<=16'd23688; ROM4[8723]<=16'd57243;
ROM1[8724]<=16'd4821; ROM2[8724]<=16'd0; ROM3[8724]<=16'd23682; ROM4[8724]<=16'd57236;
ROM1[8725]<=16'd4812; ROM2[8725]<=16'd0; ROM3[8725]<=16'd23697; ROM4[8725]<=16'd57241;
ROM1[8726]<=16'd4808; ROM2[8726]<=16'd0; ROM3[8726]<=16'd23723; ROM4[8726]<=16'd57253;
ROM1[8727]<=16'd4800; ROM2[8727]<=16'd0; ROM3[8727]<=16'd23734; ROM4[8727]<=16'd57260;
ROM1[8728]<=16'd4793; ROM2[8728]<=16'd0; ROM3[8728]<=16'd23746; ROM4[8728]<=16'd57267;
ROM1[8729]<=16'd4799; ROM2[8729]<=16'd0; ROM3[8729]<=16'd23751; ROM4[8729]<=16'd57270;
ROM1[8730]<=16'd4813; ROM2[8730]<=16'd0; ROM3[8730]<=16'd23740; ROM4[8730]<=16'd57263;
ROM1[8731]<=16'd4845; ROM2[8731]<=16'd0; ROM3[8731]<=16'd23734; ROM4[8731]<=16'd57265;
ROM1[8732]<=16'd4880; ROM2[8732]<=16'd0; ROM3[8732]<=16'd23761; ROM4[8732]<=16'd57297;
ROM1[8733]<=16'd4871; ROM2[8733]<=16'd0; ROM3[8733]<=16'd23769; ROM4[8733]<=16'd57302;
ROM1[8734]<=16'd4829; ROM2[8734]<=16'd0; ROM3[8734]<=16'd23754; ROM4[8734]<=16'd57279;
ROM1[8735]<=16'd4823; ROM2[8735]<=16'd0; ROM3[8735]<=16'd23768; ROM4[8735]<=16'd57284;
ROM1[8736]<=16'd4804; ROM2[8736]<=16'd0; ROM3[8736]<=16'd23773; ROM4[8736]<=16'd57279;
ROM1[8737]<=16'd4793; ROM2[8737]<=16'd0; ROM3[8737]<=16'd23767; ROM4[8737]<=16'd57270;
ROM1[8738]<=16'd4823; ROM2[8738]<=16'd0; ROM3[8738]<=16'd23774; ROM4[8738]<=16'd57282;
ROM1[8739]<=16'd4849; ROM2[8739]<=16'd0; ROM3[8739]<=16'd23757; ROM4[8739]<=16'd57277;
ROM1[8740]<=16'd4858; ROM2[8740]<=16'd0; ROM3[8740]<=16'd23736; ROM4[8740]<=16'd57269;
ROM1[8741]<=16'd4854; ROM2[8741]<=16'd0; ROM3[8741]<=16'd23739; ROM4[8741]<=16'd57274;
ROM1[8742]<=16'd4841; ROM2[8742]<=16'd0; ROM3[8742]<=16'd23749; ROM4[8742]<=16'd57278;
ROM1[8743]<=16'd4825; ROM2[8743]<=16'd0; ROM3[8743]<=16'd23752; ROM4[8743]<=16'd57276;
ROM1[8744]<=16'd4813; ROM2[8744]<=16'd0; ROM3[8744]<=16'd23756; ROM4[8744]<=16'd57278;
ROM1[8745]<=16'd4813; ROM2[8745]<=16'd0; ROM3[8745]<=16'd23768; ROM4[8745]<=16'd57284;
ROM1[8746]<=16'd4822; ROM2[8746]<=16'd0; ROM3[8746]<=16'd23762; ROM4[8746]<=16'd57285;
ROM1[8747]<=16'd4859; ROM2[8747]<=16'd0; ROM3[8747]<=16'd23761; ROM4[8747]<=16'd57289;
ROM1[8748]<=16'd4876; ROM2[8748]<=16'd0; ROM3[8748]<=16'd23742; ROM4[8748]<=16'd57278;
ROM1[8749]<=16'd4840; ROM2[8749]<=16'd0; ROM3[8749]<=16'd23708; ROM4[8749]<=16'd57247;
ROM1[8750]<=16'd4813; ROM2[8750]<=16'd0; ROM3[8750]<=16'd23703; ROM4[8750]<=16'd57232;
ROM1[8751]<=16'd4785; ROM2[8751]<=16'd0; ROM3[8751]<=16'd23697; ROM4[8751]<=16'd57219;
ROM1[8752]<=16'd4769; ROM2[8752]<=16'd0; ROM3[8752]<=16'd23697; ROM4[8752]<=16'd57218;
ROM1[8753]<=16'd4767; ROM2[8753]<=16'd0; ROM3[8753]<=16'd23710; ROM4[8753]<=16'd57226;
ROM1[8754]<=16'd4768; ROM2[8754]<=16'd0; ROM3[8754]<=16'd23706; ROM4[8754]<=16'd57231;
ROM1[8755]<=16'd4782; ROM2[8755]<=16'd0; ROM3[8755]<=16'd23688; ROM4[8755]<=16'd57226;
ROM1[8756]<=16'd4811; ROM2[8756]<=16'd0; ROM3[8756]<=16'd23673; ROM4[8756]<=16'd57217;
ROM1[8757]<=16'd4822; ROM2[8757]<=16'd0; ROM3[8757]<=16'd23672; ROM4[8757]<=16'd57218;
ROM1[8758]<=16'd4809; ROM2[8758]<=16'd0; ROM3[8758]<=16'd23683; ROM4[8758]<=16'd57220;
ROM1[8759]<=16'd4788; ROM2[8759]<=16'd0; ROM3[8759]<=16'd23693; ROM4[8759]<=16'd57220;
ROM1[8760]<=16'd4776; ROM2[8760]<=16'd0; ROM3[8760]<=16'd23699; ROM4[8760]<=16'd57218;
ROM1[8761]<=16'd4763; ROM2[8761]<=16'd0; ROM3[8761]<=16'd23707; ROM4[8761]<=16'd57215;
ROM1[8762]<=16'd4770; ROM2[8762]<=16'd0; ROM3[8762]<=16'd23715; ROM4[8762]<=16'd57220;
ROM1[8763]<=16'd4796; ROM2[8763]<=16'd0; ROM3[8763]<=16'd23722; ROM4[8763]<=16'd57235;
ROM1[8764]<=16'd4812; ROM2[8764]<=16'd0; ROM3[8764]<=16'd23706; ROM4[8764]<=16'd57230;
ROM1[8765]<=16'd4813; ROM2[8765]<=16'd0; ROM3[8765]<=16'd23685; ROM4[8765]<=16'd57216;
ROM1[8766]<=16'd4800; ROM2[8766]<=16'd0; ROM3[8766]<=16'd23683; ROM4[8766]<=16'd57214;
ROM1[8767]<=16'd4771; ROM2[8767]<=16'd0; ROM3[8767]<=16'd23685; ROM4[8767]<=16'd57208;
ROM1[8768]<=16'd4757; ROM2[8768]<=16'd0; ROM3[8768]<=16'd23696; ROM4[8768]<=16'd57215;
ROM1[8769]<=16'd4753; ROM2[8769]<=16'd0; ROM3[8769]<=16'd23715; ROM4[8769]<=16'd57228;
ROM1[8770]<=16'd4751; ROM2[8770]<=16'd0; ROM3[8770]<=16'd23730; ROM4[8770]<=16'd57235;
ROM1[8771]<=16'd4763; ROM2[8771]<=16'd0; ROM3[8771]<=16'd23729; ROM4[8771]<=16'd57235;
ROM1[8772]<=16'd4783; ROM2[8772]<=16'd0; ROM3[8772]<=16'd23706; ROM4[8772]<=16'd57225;
ROM1[8773]<=16'd4808; ROM2[8773]<=16'd0; ROM3[8773]<=16'd23693; ROM4[8773]<=16'd57226;
ROM1[8774]<=16'd4820; ROM2[8774]<=16'd0; ROM3[8774]<=16'd23709; ROM4[8774]<=16'd57239;
ROM1[8775]<=16'd4801; ROM2[8775]<=16'd0; ROM3[8775]<=16'd23706; ROM4[8775]<=16'd57233;
ROM1[8776]<=16'd4779; ROM2[8776]<=16'd0; ROM3[8776]<=16'd23706; ROM4[8776]<=16'd57225;
ROM1[8777]<=16'd4776; ROM2[8777]<=16'd0; ROM3[8777]<=16'd23724; ROM4[8777]<=16'd57240;
ROM1[8778]<=16'd4765; ROM2[8778]<=16'd0; ROM3[8778]<=16'd23724; ROM4[8778]<=16'd57239;
ROM1[8779]<=16'd4767; ROM2[8779]<=16'd0; ROM3[8779]<=16'd23716; ROM4[8779]<=16'd57232;
ROM1[8780]<=16'd4795; ROM2[8780]<=16'd0; ROM3[8780]<=16'd23713; ROM4[8780]<=16'd57236;
ROM1[8781]<=16'd4829; ROM2[8781]<=16'd0; ROM3[8781]<=16'd23707; ROM4[8781]<=16'd57239;
ROM1[8782]<=16'd4831; ROM2[8782]<=16'd0; ROM3[8782]<=16'd23702; ROM4[8782]<=16'd57239;
ROM1[8783]<=16'd4817; ROM2[8783]<=16'd0; ROM3[8783]<=16'd23713; ROM4[8783]<=16'd57244;
ROM1[8784]<=16'd4828; ROM2[8784]<=16'd0; ROM3[8784]<=16'd23749; ROM4[8784]<=16'd57270;
ROM1[8785]<=16'd4840; ROM2[8785]<=16'd0; ROM3[8785]<=16'd23775; ROM4[8785]<=16'd57291;
ROM1[8786]<=16'd4797; ROM2[8786]<=16'd0; ROM3[8786]<=16'd23755; ROM4[8786]<=16'd57263;
ROM1[8787]<=16'd4777; ROM2[8787]<=16'd0; ROM3[8787]<=16'd23742; ROM4[8787]<=16'd57250;
ROM1[8788]<=16'd4790; ROM2[8788]<=16'd0; ROM3[8788]<=16'd23738; ROM4[8788]<=16'd57253;
ROM1[8789]<=16'd4821; ROM2[8789]<=16'd0; ROM3[8789]<=16'd23732; ROM4[8789]<=16'd57256;
ROM1[8790]<=16'd4862; ROM2[8790]<=16'd0; ROM3[8790]<=16'd23750; ROM4[8790]<=16'd57283;
ROM1[8791]<=16'd4860; ROM2[8791]<=16'd0; ROM3[8791]<=16'd23767; ROM4[8791]<=16'd57294;
ROM1[8792]<=16'd4834; ROM2[8792]<=16'd0; ROM3[8792]<=16'd23770; ROM4[8792]<=16'd57290;
ROM1[8793]<=16'd4808; ROM2[8793]<=16'd0; ROM3[8793]<=16'd23767; ROM4[8793]<=16'd57282;
ROM1[8794]<=16'd4782; ROM2[8794]<=16'd0; ROM3[8794]<=16'd23765; ROM4[8794]<=16'd57274;
ROM1[8795]<=16'd4774; ROM2[8795]<=16'd0; ROM3[8795]<=16'd23770; ROM4[8795]<=16'd57274;
ROM1[8796]<=16'd4786; ROM2[8796]<=16'd0; ROM3[8796]<=16'd23772; ROM4[8796]<=16'd57275;
ROM1[8797]<=16'd4815; ROM2[8797]<=16'd0; ROM3[8797]<=16'd23759; ROM4[8797]<=16'd57276;
ROM1[8798]<=16'd4844; ROM2[8798]<=16'd0; ROM3[8798]<=16'd23747; ROM4[8798]<=16'd57276;
ROM1[8799]<=16'd4851; ROM2[8799]<=16'd0; ROM3[8799]<=16'd23751; ROM4[8799]<=16'd57278;
ROM1[8800]<=16'd4844; ROM2[8800]<=16'd0; ROM3[8800]<=16'd23759; ROM4[8800]<=16'd57283;
ROM1[8801]<=16'd4814; ROM2[8801]<=16'd0; ROM3[8801]<=16'd23752; ROM4[8801]<=16'd57270;
ROM1[8802]<=16'd4791; ROM2[8802]<=16'd0; ROM3[8802]<=16'd23743; ROM4[8802]<=16'd57256;
ROM1[8803]<=16'd4784; ROM2[8803]<=16'd0; ROM3[8803]<=16'd23752; ROM4[8803]<=16'd57262;
ROM1[8804]<=16'd4782; ROM2[8804]<=16'd0; ROM3[8804]<=16'd23745; ROM4[8804]<=16'd57253;
ROM1[8805]<=16'd4801; ROM2[8805]<=16'd0; ROM3[8805]<=16'd23735; ROM4[8805]<=16'd57245;
ROM1[8806]<=16'd4840; ROM2[8806]<=16'd0; ROM3[8806]<=16'd23734; ROM4[8806]<=16'd57256;
ROM1[8807]<=16'd4845; ROM2[8807]<=16'd0; ROM3[8807]<=16'd23732; ROM4[8807]<=16'd57258;
ROM1[8808]<=16'd4833; ROM2[8808]<=16'd0; ROM3[8808]<=16'd23741; ROM4[8808]<=16'd57266;
ROM1[8809]<=16'd4824; ROM2[8809]<=16'd0; ROM3[8809]<=16'd23761; ROM4[8809]<=16'd57273;
ROM1[8810]<=16'd4813; ROM2[8810]<=16'd0; ROM3[8810]<=16'd23774; ROM4[8810]<=16'd57279;
ROM1[8811]<=16'd4794; ROM2[8811]<=16'd0; ROM3[8811]<=16'd23778; ROM4[8811]<=16'd57280;
ROM1[8812]<=16'd4795; ROM2[8812]<=16'd0; ROM3[8812]<=16'd23785; ROM4[8812]<=16'd57287;
ROM1[8813]<=16'd4821; ROM2[8813]<=16'd0; ROM3[8813]<=16'd23787; ROM4[8813]<=16'd57297;
ROM1[8814]<=16'd4854; ROM2[8814]<=16'd0; ROM3[8814]<=16'd23777; ROM4[8814]<=16'd57301;
ROM1[8815]<=16'd4877; ROM2[8815]<=16'd0; ROM3[8815]<=16'd23776; ROM4[8815]<=16'd57307;
ROM1[8816]<=16'd4851; ROM2[8816]<=16'd0; ROM3[8816]<=16'd23769; ROM4[8816]<=16'd57293;
ROM1[8817]<=16'd4820; ROM2[8817]<=16'd0; ROM3[8817]<=16'd23762; ROM4[8817]<=16'd57281;
ROM1[8818]<=16'd4799; ROM2[8818]<=16'd0; ROM3[8818]<=16'd23759; ROM4[8818]<=16'd57275;
ROM1[8819]<=16'd4769; ROM2[8819]<=16'd0; ROM3[8819]<=16'd23746; ROM4[8819]<=16'd57254;
ROM1[8820]<=16'd4761; ROM2[8820]<=16'd0; ROM3[8820]<=16'd23740; ROM4[8820]<=16'd57249;
ROM1[8821]<=16'd4771; ROM2[8821]<=16'd0; ROM3[8821]<=16'd23733; ROM4[8821]<=16'd57247;
ROM1[8822]<=16'd4794; ROM2[8822]<=16'd0; ROM3[8822]<=16'd23719; ROM4[8822]<=16'd57239;
ROM1[8823]<=16'd4817; ROM2[8823]<=16'd0; ROM3[8823]<=16'd23701; ROM4[8823]<=16'd57236;
ROM1[8824]<=16'd4808; ROM2[8824]<=16'd0; ROM3[8824]<=16'd23691; ROM4[8824]<=16'd57226;
ROM1[8825]<=16'd4792; ROM2[8825]<=16'd0; ROM3[8825]<=16'd23695; ROM4[8825]<=16'd57225;
ROM1[8826]<=16'd4780; ROM2[8826]<=16'd0; ROM3[8826]<=16'd23704; ROM4[8826]<=16'd57228;
ROM1[8827]<=16'd4775; ROM2[8827]<=16'd0; ROM3[8827]<=16'd23715; ROM4[8827]<=16'd57236;
ROM1[8828]<=16'd4771; ROM2[8828]<=16'd0; ROM3[8828]<=16'd23726; ROM4[8828]<=16'd57246;
ROM1[8829]<=16'd4779; ROM2[8829]<=16'd0; ROM3[8829]<=16'd23736; ROM4[8829]<=16'd57253;
ROM1[8830]<=16'd4796; ROM2[8830]<=16'd0; ROM3[8830]<=16'd23724; ROM4[8830]<=16'd57246;
ROM1[8831]<=16'd4812; ROM2[8831]<=16'd0; ROM3[8831]<=16'd23699; ROM4[8831]<=16'd57233;
ROM1[8832]<=16'd4813; ROM2[8832]<=16'd0; ROM3[8832]<=16'd23699; ROM4[8832]<=16'd57234;
ROM1[8833]<=16'd4798; ROM2[8833]<=16'd0; ROM3[8833]<=16'd23701; ROM4[8833]<=16'd57234;
ROM1[8834]<=16'd4772; ROM2[8834]<=16'd0; ROM3[8834]<=16'd23695; ROM4[8834]<=16'd57226;
ROM1[8835]<=16'd4762; ROM2[8835]<=16'd0; ROM3[8835]<=16'd23712; ROM4[8835]<=16'd57227;
ROM1[8836]<=16'd4756; ROM2[8836]<=16'd0; ROM3[8836]<=16'd23732; ROM4[8836]<=16'd57234;
ROM1[8837]<=16'd4746; ROM2[8837]<=16'd0; ROM3[8837]<=16'd23731; ROM4[8837]<=16'd57233;
ROM1[8838]<=16'd4770; ROM2[8838]<=16'd0; ROM3[8838]<=16'd23739; ROM4[8838]<=16'd57246;
ROM1[8839]<=16'd4812; ROM2[8839]<=16'd0; ROM3[8839]<=16'd23734; ROM4[8839]<=16'd57252;
ROM1[8840]<=16'd4824; ROM2[8840]<=16'd0; ROM3[8840]<=16'd23723; ROM4[8840]<=16'd57244;
ROM1[8841]<=16'd4823; ROM2[8841]<=16'd0; ROM3[8841]<=16'd23741; ROM4[8841]<=16'd57254;
ROM1[8842]<=16'd4823; ROM2[8842]<=16'd0; ROM3[8842]<=16'd23769; ROM4[8842]<=16'd57276;
ROM1[8843]<=16'd4805; ROM2[8843]<=16'd0; ROM3[8843]<=16'd23773; ROM4[8843]<=16'd57273;
ROM1[8844]<=16'd4782; ROM2[8844]<=16'd0; ROM3[8844]<=16'd23770; ROM4[8844]<=16'd57268;
ROM1[8845]<=16'd4773; ROM2[8845]<=16'd0; ROM3[8845]<=16'd23766; ROM4[8845]<=16'd57263;
ROM1[8846]<=16'd4779; ROM2[8846]<=16'd0; ROM3[8846]<=16'd23755; ROM4[8846]<=16'd57256;
ROM1[8847]<=16'd4808; ROM2[8847]<=16'd0; ROM3[8847]<=16'd23743; ROM4[8847]<=16'd57254;
ROM1[8848]<=16'd4835; ROM2[8848]<=16'd0; ROM3[8848]<=16'd23731; ROM4[8848]<=16'd57254;
ROM1[8849]<=16'd4833; ROM2[8849]<=16'd0; ROM3[8849]<=16'd23731; ROM4[8849]<=16'd57257;
ROM1[8850]<=16'd4825; ROM2[8850]<=16'd0; ROM3[8850]<=16'd23747; ROM4[8850]<=16'd57270;
ROM1[8851]<=16'd4824; ROM2[8851]<=16'd0; ROM3[8851]<=16'd23768; ROM4[8851]<=16'd57286;
ROM1[8852]<=16'd4804; ROM2[8852]<=16'd0; ROM3[8852]<=16'd23761; ROM4[8852]<=16'd57278;
ROM1[8853]<=16'd4782; ROM2[8853]<=16'd0; ROM3[8853]<=16'd23755; ROM4[8853]<=16'd57267;
ROM1[8854]<=16'd4773; ROM2[8854]<=16'd0; ROM3[8854]<=16'd23743; ROM4[8854]<=16'd57252;
ROM1[8855]<=16'd4785; ROM2[8855]<=16'd0; ROM3[8855]<=16'd23726; ROM4[8855]<=16'd57247;
ROM1[8856]<=16'd4824; ROM2[8856]<=16'd0; ROM3[8856]<=16'd23719; ROM4[8856]<=16'd57257;
ROM1[8857]<=16'd4832; ROM2[8857]<=16'd0; ROM3[8857]<=16'd23705; ROM4[8857]<=16'd57246;
ROM1[8858]<=16'd4815; ROM2[8858]<=16'd0; ROM3[8858]<=16'd23701; ROM4[8858]<=16'd57237;
ROM1[8859]<=16'd4805; ROM2[8859]<=16'd0; ROM3[8859]<=16'd23715; ROM4[8859]<=16'd57239;
ROM1[8860]<=16'd4793; ROM2[8860]<=16'd0; ROM3[8860]<=16'd23726; ROM4[8860]<=16'd57239;
ROM1[8861]<=16'd4769; ROM2[8861]<=16'd0; ROM3[8861]<=16'd23735; ROM4[8861]<=16'd57239;
ROM1[8862]<=16'd4764; ROM2[8862]<=16'd0; ROM3[8862]<=16'd23741; ROM4[8862]<=16'd57245;
ROM1[8863]<=16'd4777; ROM2[8863]<=16'd0; ROM3[8863]<=16'd23727; ROM4[8863]<=16'd57240;
ROM1[8864]<=16'd4807; ROM2[8864]<=16'd0; ROM3[8864]<=16'd23717; ROM4[8864]<=16'd57237;
ROM1[8865]<=16'd4824; ROM2[8865]<=16'd0; ROM3[8865]<=16'd23706; ROM4[8865]<=16'd57235;
ROM1[8866]<=16'd4809; ROM2[8866]<=16'd0; ROM3[8866]<=16'd23702; ROM4[8866]<=16'd57229;
ROM1[8867]<=16'd4796; ROM2[8867]<=16'd0; ROM3[8867]<=16'd23722; ROM4[8867]<=16'd57238;
ROM1[8868]<=16'd4807; ROM2[8868]<=16'd0; ROM3[8868]<=16'd23752; ROM4[8868]<=16'd57264;
ROM1[8869]<=16'd4793; ROM2[8869]<=16'd0; ROM3[8869]<=16'd23756; ROM4[8869]<=16'd57266;
ROM1[8870]<=16'd4767; ROM2[8870]<=16'd0; ROM3[8870]<=16'd23736; ROM4[8870]<=16'd57245;
ROM1[8871]<=16'd4762; ROM2[8871]<=16'd0; ROM3[8871]<=16'd23715; ROM4[8871]<=16'd57232;
ROM1[8872]<=16'd4778; ROM2[8872]<=16'd0; ROM3[8872]<=16'd23699; ROM4[8872]<=16'd57226;
ROM1[8873]<=16'd4807; ROM2[8873]<=16'd0; ROM3[8873]<=16'd23691; ROM4[8873]<=16'd57228;
ROM1[8874]<=16'd4823; ROM2[8874]<=16'd0; ROM3[8874]<=16'd23707; ROM4[8874]<=16'd57243;
ROM1[8875]<=16'd4818; ROM2[8875]<=16'd0; ROM3[8875]<=16'd23723; ROM4[8875]<=16'd57251;
ROM1[8876]<=16'd4782; ROM2[8876]<=16'd0; ROM3[8876]<=16'd23712; ROM4[8876]<=16'd57235;
ROM1[8877]<=16'd4766; ROM2[8877]<=16'd0; ROM3[8877]<=16'd23716; ROM4[8877]<=16'd57233;
ROM1[8878]<=16'd4756; ROM2[8878]<=16'd0; ROM3[8878]<=16'd23726; ROM4[8878]<=16'd57234;
ROM1[8879]<=16'd4758; ROM2[8879]<=16'd0; ROM3[8879]<=16'd23718; ROM4[8879]<=16'd57227;
ROM1[8880]<=16'd4783; ROM2[8880]<=16'd0; ROM3[8880]<=16'd23704; ROM4[8880]<=16'd57225;
ROM1[8881]<=16'd4814; ROM2[8881]<=16'd0; ROM3[8881]<=16'd23698; ROM4[8881]<=16'd57229;
ROM1[8882]<=16'd4825; ROM2[8882]<=16'd0; ROM3[8882]<=16'd23704; ROM4[8882]<=16'd57234;
ROM1[8883]<=16'd4808; ROM2[8883]<=16'd0; ROM3[8883]<=16'd23710; ROM4[8883]<=16'd57237;
ROM1[8884]<=16'd4786; ROM2[8884]<=16'd0; ROM3[8884]<=16'd23718; ROM4[8884]<=16'd57236;
ROM1[8885]<=16'd4783; ROM2[8885]<=16'd0; ROM3[8885]<=16'd23727; ROM4[8885]<=16'd57243;
ROM1[8886]<=16'd4790; ROM2[8886]<=16'd0; ROM3[8886]<=16'd23749; ROM4[8886]<=16'd57262;
ROM1[8887]<=16'd4787; ROM2[8887]<=16'd0; ROM3[8887]<=16'd23747; ROM4[8887]<=16'd57259;
ROM1[8888]<=16'd4790; ROM2[8888]<=16'd0; ROM3[8888]<=16'd23723; ROM4[8888]<=16'd57243;
ROM1[8889]<=16'd4815; ROM2[8889]<=16'd0; ROM3[8889]<=16'd23706; ROM4[8889]<=16'd57234;
ROM1[8890]<=16'd4818; ROM2[8890]<=16'd0; ROM3[8890]<=16'd23685; ROM4[8890]<=16'd57220;
ROM1[8891]<=16'd4806; ROM2[8891]<=16'd0; ROM3[8891]<=16'd23685; ROM4[8891]<=16'd57219;
ROM1[8892]<=16'd4808; ROM2[8892]<=16'd0; ROM3[8892]<=16'd23711; ROM4[8892]<=16'd57241;
ROM1[8893]<=16'd4812; ROM2[8893]<=16'd0; ROM3[8893]<=16'd23737; ROM4[8893]<=16'd57260;
ROM1[8894]<=16'd4795; ROM2[8894]<=16'd0; ROM3[8894]<=16'd23740; ROM4[8894]<=16'd57259;
ROM1[8895]<=16'd4792; ROM2[8895]<=16'd0; ROM3[8895]<=16'd23748; ROM4[8895]<=16'd57261;
ROM1[8896]<=16'd4813; ROM2[8896]<=16'd0; ROM3[8896]<=16'd23757; ROM4[8896]<=16'd57271;
ROM1[8897]<=16'd4825; ROM2[8897]<=16'd0; ROM3[8897]<=16'd23732; ROM4[8897]<=16'd57255;
ROM1[8898]<=16'd4846; ROM2[8898]<=16'd0; ROM3[8898]<=16'd23721; ROM4[8898]<=16'd57253;
ROM1[8899]<=16'd4842; ROM2[8899]<=16'd0; ROM3[8899]<=16'd23725; ROM4[8899]<=16'd57257;
ROM1[8900]<=16'd4845; ROM2[8900]<=16'd0; ROM3[8900]<=16'd23744; ROM4[8900]<=16'd57269;
ROM1[8901]<=16'd4850; ROM2[8901]<=16'd0; ROM3[8901]<=16'd23765; ROM4[8901]<=16'd57284;
ROM1[8902]<=16'd4805; ROM2[8902]<=16'd0; ROM3[8902]<=16'd23737; ROM4[8902]<=16'd57254;
ROM1[8903]<=16'd4778; ROM2[8903]<=16'd0; ROM3[8903]<=16'd23730; ROM4[8903]<=16'd57236;
ROM1[8904]<=16'd4774; ROM2[8904]<=16'd0; ROM3[8904]<=16'd23721; ROM4[8904]<=16'd57226;
ROM1[8905]<=16'd4790; ROM2[8905]<=16'd0; ROM3[8905]<=16'd23709; ROM4[8905]<=16'd57223;
ROM1[8906]<=16'd4849; ROM2[8906]<=16'd0; ROM3[8906]<=16'd23724; ROM4[8906]<=16'd57249;
ROM1[8907]<=16'd4862; ROM2[8907]<=16'd0; ROM3[8907]<=16'd23726; ROM4[8907]<=16'd57257;
ROM1[8908]<=16'd4823; ROM2[8908]<=16'd0; ROM3[8908]<=16'd23707; ROM4[8908]<=16'd57234;
ROM1[8909]<=16'd4795; ROM2[8909]<=16'd0; ROM3[8909]<=16'd23705; ROM4[8909]<=16'd57223;
ROM1[8910]<=16'd4790; ROM2[8910]<=16'd0; ROM3[8910]<=16'd23715; ROM4[8910]<=16'd57231;
ROM1[8911]<=16'd4777; ROM2[8911]<=16'd0; ROM3[8911]<=16'd23720; ROM4[8911]<=16'd57235;
ROM1[8912]<=16'd4770; ROM2[8912]<=16'd0; ROM3[8912]<=16'd23714; ROM4[8912]<=16'd57231;
ROM1[8913]<=16'd4776; ROM2[8913]<=16'd0; ROM3[8913]<=16'd23698; ROM4[8913]<=16'd57219;
ROM1[8914]<=16'd4797; ROM2[8914]<=16'd0; ROM3[8914]<=16'd23679; ROM4[8914]<=16'd57211;
ROM1[8915]<=16'd4818; ROM2[8915]<=16'd0; ROM3[8915]<=16'd23674; ROM4[8915]<=16'd57213;
ROM1[8916]<=16'd4810; ROM2[8916]<=16'd0; ROM3[8916]<=16'd23683; ROM4[8916]<=16'd57220;
ROM1[8917]<=16'd4781; ROM2[8917]<=16'd0; ROM3[8917]<=16'd23684; ROM4[8917]<=16'd57214;
ROM1[8918]<=16'd4763; ROM2[8918]<=16'd0; ROM3[8918]<=16'd23686; ROM4[8918]<=16'd57205;
ROM1[8919]<=16'd4743; ROM2[8919]<=16'd0; ROM3[8919]<=16'd23686; ROM4[8919]<=16'd57199;
ROM1[8920]<=16'd4749; ROM2[8920]<=16'd0; ROM3[8920]<=16'd23699; ROM4[8920]<=16'd57206;
ROM1[8921]<=16'd4774; ROM2[8921]<=16'd0; ROM3[8921]<=16'd23707; ROM4[8921]<=16'd57219;
ROM1[8922]<=16'd4791; ROM2[8922]<=16'd0; ROM3[8922]<=16'd23686; ROM4[8922]<=16'd57208;
ROM1[8923]<=16'd4802; ROM2[8923]<=16'd0; ROM3[8923]<=16'd23663; ROM4[8923]<=16'd57196;
ROM1[8924]<=16'd4795; ROM2[8924]<=16'd0; ROM3[8924]<=16'd23656; ROM4[8924]<=16'd57194;
ROM1[8925]<=16'd4779; ROM2[8925]<=16'd0; ROM3[8925]<=16'd23662; ROM4[8925]<=16'd57195;
ROM1[8926]<=16'd4766; ROM2[8926]<=16'd0; ROM3[8926]<=16'd23671; ROM4[8926]<=16'd57196;
ROM1[8927]<=16'd4762; ROM2[8927]<=16'd0; ROM3[8927]<=16'd23679; ROM4[8927]<=16'd57203;
ROM1[8928]<=16'd4751; ROM2[8928]<=16'd0; ROM3[8928]<=16'd23683; ROM4[8928]<=16'd57205;
ROM1[8929]<=16'd4753; ROM2[8929]<=16'd0; ROM3[8929]<=16'd23683; ROM4[8929]<=16'd57205;
ROM1[8930]<=16'd4779; ROM2[8930]<=16'd0; ROM3[8930]<=16'd23680; ROM4[8930]<=16'd57208;
ROM1[8931]<=16'd4816; ROM2[8931]<=16'd0; ROM3[8931]<=16'd23678; ROM4[8931]<=16'd57220;
ROM1[8932]<=16'd4829; ROM2[8932]<=16'd0; ROM3[8932]<=16'd23686; ROM4[8932]<=16'd57229;
ROM1[8933]<=16'd4832; ROM2[8933]<=16'd0; ROM3[8933]<=16'd23704; ROM4[8933]<=16'd57240;
ROM1[8934]<=16'd4816; ROM2[8934]<=16'd0; ROM3[8934]<=16'd23715; ROM4[8934]<=16'd57247;
ROM1[8935]<=16'd4795; ROM2[8935]<=16'd0; ROM3[8935]<=16'd23720; ROM4[8935]<=16'd57244;
ROM1[8936]<=16'd4795; ROM2[8936]<=16'd0; ROM3[8936]<=16'd23743; ROM4[8936]<=16'd57256;
ROM1[8937]<=16'd4789; ROM2[8937]<=16'd0; ROM3[8937]<=16'd23744; ROM4[8937]<=16'd57252;
ROM1[8938]<=16'd4784; ROM2[8938]<=16'd0; ROM3[8938]<=16'd23720; ROM4[8938]<=16'd57231;
ROM1[8939]<=16'd4817; ROM2[8939]<=16'd0; ROM3[8939]<=16'd23703; ROM4[8939]<=16'd57226;
ROM1[8940]<=16'd4823; ROM2[8940]<=16'd0; ROM3[8940]<=16'd23692; ROM4[8940]<=16'd57218;
ROM1[8941]<=16'd4801; ROM2[8941]<=16'd0; ROM3[8941]<=16'd23689; ROM4[8941]<=16'd57211;
ROM1[8942]<=16'd4800; ROM2[8942]<=16'd0; ROM3[8942]<=16'd23711; ROM4[8942]<=16'd57228;
ROM1[8943]<=16'd4787; ROM2[8943]<=16'd0; ROM3[8943]<=16'd23723; ROM4[8943]<=16'd57231;
ROM1[8944]<=16'd4764; ROM2[8944]<=16'd0; ROM3[8944]<=16'd23719; ROM4[8944]<=16'd57226;
ROM1[8945]<=16'd4764; ROM2[8945]<=16'd0; ROM3[8945]<=16'd23723; ROM4[8945]<=16'd57229;
ROM1[8946]<=16'd4785; ROM2[8946]<=16'd0; ROM3[8946]<=16'd23728; ROM4[8946]<=16'd57238;
ROM1[8947]<=16'd4812; ROM2[8947]<=16'd0; ROM3[8947]<=16'd23722; ROM4[8947]<=16'd57242;
ROM1[8948]<=16'd4832; ROM2[8948]<=16'd0; ROM3[8948]<=16'd23706; ROM4[8948]<=16'd57238;
ROM1[8949]<=16'd4829; ROM2[8949]<=16'd0; ROM3[8949]<=16'd23709; ROM4[8949]<=16'd57239;
ROM1[8950]<=16'd4813; ROM2[8950]<=16'd0; ROM3[8950]<=16'd23719; ROM4[8950]<=16'd57239;
ROM1[8951]<=16'd4799; ROM2[8951]<=16'd0; ROM3[8951]<=16'd23730; ROM4[8951]<=16'd57242;
ROM1[8952]<=16'd4795; ROM2[8952]<=16'd0; ROM3[8952]<=16'd23744; ROM4[8952]<=16'd57255;
ROM1[8953]<=16'd4810; ROM2[8953]<=16'd0; ROM3[8953]<=16'd23772; ROM4[8953]<=16'd57280;
ROM1[8954]<=16'd4836; ROM2[8954]<=16'd0; ROM3[8954]<=16'd23790; ROM4[8954]<=16'd57302;
ROM1[8955]<=16'd4838; ROM2[8955]<=16'd0; ROM3[8955]<=16'd23754; ROM4[8955]<=16'd57278;
ROM1[8956]<=16'd4842; ROM2[8956]<=16'd0; ROM3[8956]<=16'd23713; ROM4[8956]<=16'd57245;
ROM1[8957]<=16'd4836; ROM2[8957]<=16'd0; ROM3[8957]<=16'd23701; ROM4[8957]<=16'd57235;
ROM1[8958]<=16'd4817; ROM2[8958]<=16'd0; ROM3[8958]<=16'd23699; ROM4[8958]<=16'd57230;
ROM1[8959]<=16'd4809; ROM2[8959]<=16'd0; ROM3[8959]<=16'd23718; ROM4[8959]<=16'd57241;
ROM1[8960]<=16'd4809; ROM2[8960]<=16'd0; ROM3[8960]<=16'd23740; ROM4[8960]<=16'd57257;
ROM1[8961]<=16'd4784; ROM2[8961]<=16'd0; ROM3[8961]<=16'd23737; ROM4[8961]<=16'd57248;
ROM1[8962]<=16'd4771; ROM2[8962]<=16'd0; ROM3[8962]<=16'd23728; ROM4[8962]<=16'd57243;
ROM1[8963]<=16'd4800; ROM2[8963]<=16'd0; ROM3[8963]<=16'd23730; ROM4[8963]<=16'd57252;
ROM1[8964]<=16'd4832; ROM2[8964]<=16'd0; ROM3[8964]<=16'd23719; ROM4[8964]<=16'd57249;
ROM1[8965]<=16'd4844; ROM2[8965]<=16'd0; ROM3[8965]<=16'd23708; ROM4[8965]<=16'd57251;
ROM1[8966]<=16'd4836; ROM2[8966]<=16'd0; ROM3[8966]<=16'd23719; ROM4[8966]<=16'd57257;
ROM1[8967]<=16'd4821; ROM2[8967]<=16'd0; ROM3[8967]<=16'd23734; ROM4[8967]<=16'd57263;
ROM1[8968]<=16'd4798; ROM2[8968]<=16'd0; ROM3[8968]<=16'd23733; ROM4[8968]<=16'd57255;
ROM1[8969]<=16'd4778; ROM2[8969]<=16'd0; ROM3[8969]<=16'd23735; ROM4[8969]<=16'd57249;
ROM1[8970]<=16'd4771; ROM2[8970]<=16'd0; ROM3[8970]<=16'd23740; ROM4[8970]<=16'd57252;
ROM1[8971]<=16'd4763; ROM2[8971]<=16'd0; ROM3[8971]<=16'd23723; ROM4[8971]<=16'd57235;
ROM1[8972]<=16'd4788; ROM2[8972]<=16'd0; ROM3[8972]<=16'd23711; ROM4[8972]<=16'd57232;
ROM1[8973]<=16'd4816; ROM2[8973]<=16'd0; ROM3[8973]<=16'd23701; ROM4[8973]<=16'd57232;
ROM1[8974]<=16'd4811; ROM2[8974]<=16'd0; ROM3[8974]<=16'd23698; ROM4[8974]<=16'd57227;
ROM1[8975]<=16'd4805; ROM2[8975]<=16'd0; ROM3[8975]<=16'd23716; ROM4[8975]<=16'd57236;
ROM1[8976]<=16'd4806; ROM2[8976]<=16'd0; ROM3[8976]<=16'd23743; ROM4[8976]<=16'd57253;
ROM1[8977]<=16'd4801; ROM2[8977]<=16'd0; ROM3[8977]<=16'd23757; ROM4[8977]<=16'd57263;
ROM1[8978]<=16'd4771; ROM2[8978]<=16'd0; ROM3[8978]<=16'd23740; ROM4[8978]<=16'd57242;
ROM1[8979]<=16'd4772; ROM2[8979]<=16'd0; ROM3[8979]<=16'd23735; ROM4[8979]<=16'd57236;
ROM1[8980]<=16'd4798; ROM2[8980]<=16'd0; ROM3[8980]<=16'd23731; ROM4[8980]<=16'd57241;
ROM1[8981]<=16'd4817; ROM2[8981]<=16'd0; ROM3[8981]<=16'd23710; ROM4[8981]<=16'd57229;
ROM1[8982]<=16'd4826; ROM2[8982]<=16'd0; ROM3[8982]<=16'd23710; ROM4[8982]<=16'd57231;
ROM1[8983]<=16'd4824; ROM2[8983]<=16'd0; ROM3[8983]<=16'd23729; ROM4[8983]<=16'd57247;
ROM1[8984]<=16'd4821; ROM2[8984]<=16'd0; ROM3[8984]<=16'd23748; ROM4[8984]<=16'd57260;
ROM1[8985]<=16'd4799; ROM2[8985]<=16'd0; ROM3[8985]<=16'd23743; ROM4[8985]<=16'd57249;
ROM1[8986]<=16'd4769; ROM2[8986]<=16'd0; ROM3[8986]<=16'd23733; ROM4[8986]<=16'd57237;
ROM1[8987]<=16'd4760; ROM2[8987]<=16'd0; ROM3[8987]<=16'd23727; ROM4[8987]<=16'd57232;
ROM1[8988]<=16'd4766; ROM2[8988]<=16'd0; ROM3[8988]<=16'd23710; ROM4[8988]<=16'd57223;
ROM1[8989]<=16'd4798; ROM2[8989]<=16'd0; ROM3[8989]<=16'd23700; ROM4[8989]<=16'd57227;
ROM1[8990]<=16'd4824; ROM2[8990]<=16'd0; ROM3[8990]<=16'd23697; ROM4[8990]<=16'd57233;
ROM1[8991]<=16'd4820; ROM2[8991]<=16'd0; ROM3[8991]<=16'd23698; ROM4[8991]<=16'd57234;
ROM1[8992]<=16'd4798; ROM2[8992]<=16'd0; ROM3[8992]<=16'd23698; ROM4[8992]<=16'd57231;
ROM1[8993]<=16'd4796; ROM2[8993]<=16'd0; ROM3[8993]<=16'd23717; ROM4[8993]<=16'd57241;
ROM1[8994]<=16'd4798; ROM2[8994]<=16'd0; ROM3[8994]<=16'd23746; ROM4[8994]<=16'd57262;
ROM1[8995]<=16'd4795; ROM2[8995]<=16'd0; ROM3[8995]<=16'd23755; ROM4[8995]<=16'd57268;
ROM1[8996]<=16'd4798; ROM2[8996]<=16'd0; ROM3[8996]<=16'd23748; ROM4[8996]<=16'd57259;
ROM1[8997]<=16'd4816; ROM2[8997]<=16'd0; ROM3[8997]<=16'd23726; ROM4[8997]<=16'd57248;
ROM1[8998]<=16'd4835; ROM2[8998]<=16'd0; ROM3[8998]<=16'd23708; ROM4[8998]<=16'd57239;
ROM1[8999]<=16'd4841; ROM2[8999]<=16'd0; ROM3[8999]<=16'd23722; ROM4[8999]<=16'd57254;
ROM1[9000]<=16'd4834; ROM2[9000]<=16'd0; ROM3[9000]<=16'd23736; ROM4[9000]<=16'd57266;
ROM1[9001]<=16'd4801; ROM2[9001]<=16'd0; ROM3[9001]<=16'd23725; ROM4[9001]<=16'd57248;
ROM1[9002]<=16'd4778; ROM2[9002]<=16'd0; ROM3[9002]<=16'd23725; ROM4[9002]<=16'd57241;
ROM1[9003]<=16'd4773; ROM2[9003]<=16'd0; ROM3[9003]<=16'd23733; ROM4[9003]<=16'd57248;
ROM1[9004]<=16'd4783; ROM2[9004]<=16'd0; ROM3[9004]<=16'd23734; ROM4[9004]<=16'd57250;
ROM1[9005]<=16'd4802; ROM2[9005]<=16'd0; ROM3[9005]<=16'd23724; ROM4[9005]<=16'd57243;
ROM1[9006]<=16'd4827; ROM2[9006]<=16'd0; ROM3[9006]<=16'd23708; ROM4[9006]<=16'd57240;
ROM1[9007]<=16'd4823; ROM2[9007]<=16'd0; ROM3[9007]<=16'd23694; ROM4[9007]<=16'd57228;
ROM1[9008]<=16'd4806; ROM2[9008]<=16'd0; ROM3[9008]<=16'd23696; ROM4[9008]<=16'd57223;
ROM1[9009]<=16'd4803; ROM2[9009]<=16'd0; ROM3[9009]<=16'd23725; ROM4[9009]<=16'd57243;
ROM1[9010]<=16'd4800; ROM2[9010]<=16'd0; ROM3[9010]<=16'd23741; ROM4[9010]<=16'd57254;
ROM1[9011]<=16'd4775; ROM2[9011]<=16'd0; ROM3[9011]<=16'd23744; ROM4[9011]<=16'd57245;
ROM1[9012]<=16'd4763; ROM2[9012]<=16'd0; ROM3[9012]<=16'd23743; ROM4[9012]<=16'd57238;
ROM1[9013]<=16'd4788; ROM2[9013]<=16'd0; ROM3[9013]<=16'd23742; ROM4[9013]<=16'd57242;
ROM1[9014]<=16'd4836; ROM2[9014]<=16'd0; ROM3[9014]<=16'd23753; ROM4[9014]<=16'd57257;
ROM1[9015]<=16'd4856; ROM2[9015]<=16'd0; ROM3[9015]<=16'd23748; ROM4[9015]<=16'd57260;
ROM1[9016]<=16'd4838; ROM2[9016]<=16'd0; ROM3[9016]<=16'd23743; ROM4[9016]<=16'd57257;
ROM1[9017]<=16'd4820; ROM2[9017]<=16'd0; ROM3[9017]<=16'd23751; ROM4[9017]<=16'd57265;
ROM1[9018]<=16'd4800; ROM2[9018]<=16'd0; ROM3[9018]<=16'd23753; ROM4[9018]<=16'd57265;
ROM1[9019]<=16'd4775; ROM2[9019]<=16'd0; ROM3[9019]<=16'd23750; ROM4[9019]<=16'd57256;
ROM1[9020]<=16'd4763; ROM2[9020]<=16'd0; ROM3[9020]<=16'd23745; ROM4[9020]<=16'd57252;
ROM1[9021]<=16'd4764; ROM2[9021]<=16'd0; ROM3[9021]<=16'd23730; ROM4[9021]<=16'd57240;
ROM1[9022]<=16'd4786; ROM2[9022]<=16'd0; ROM3[9022]<=16'd23709; ROM4[9022]<=16'd57228;
ROM1[9023]<=16'd4806; ROM2[9023]<=16'd0; ROM3[9023]<=16'd23692; ROM4[9023]<=16'd57227;
ROM1[9024]<=16'd4802; ROM2[9024]<=16'd0; ROM3[9024]<=16'd23695; ROM4[9024]<=16'd57230;
ROM1[9025]<=16'd4793; ROM2[9025]<=16'd0; ROM3[9025]<=16'd23708; ROM4[9025]<=16'd57238;
ROM1[9026]<=16'd4781; ROM2[9026]<=16'd0; ROM3[9026]<=16'd23715; ROM4[9026]<=16'd57241;
ROM1[9027]<=16'd4768; ROM2[9027]<=16'd0; ROM3[9027]<=16'd23717; ROM4[9027]<=16'd57237;
ROM1[9028]<=16'd4761; ROM2[9028]<=16'd0; ROM3[9028]<=16'd23719; ROM4[9028]<=16'd57236;
ROM1[9029]<=16'd4775; ROM2[9029]<=16'd0; ROM3[9029]<=16'd23726; ROM4[9029]<=16'd57246;
ROM1[9030]<=16'd4813; ROM2[9030]<=16'd0; ROM3[9030]<=16'd23734; ROM4[9030]<=16'd57261;
ROM1[9031]<=16'd4853; ROM2[9031]<=16'd0; ROM3[9031]<=16'd23731; ROM4[9031]<=16'd57269;
ROM1[9032]<=16'd4844; ROM2[9032]<=16'd0; ROM3[9032]<=16'd23713; ROM4[9032]<=16'd57255;
ROM1[9033]<=16'd4813; ROM2[9033]<=16'd0; ROM3[9033]<=16'd23700; ROM4[9033]<=16'd57234;
ROM1[9034]<=16'd4789; ROM2[9034]<=16'd0; ROM3[9034]<=16'd23701; ROM4[9034]<=16'd57223;
ROM1[9035]<=16'd4785; ROM2[9035]<=16'd0; ROM3[9035]<=16'd23718; ROM4[9035]<=16'd57232;
ROM1[9036]<=16'd4792; ROM2[9036]<=16'd0; ROM3[9036]<=16'd23747; ROM4[9036]<=16'd57253;
ROM1[9037]<=16'd4778; ROM2[9037]<=16'd0; ROM3[9037]<=16'd23732; ROM4[9037]<=16'd57238;
ROM1[9038]<=16'd4769; ROM2[9038]<=16'd0; ROM3[9038]<=16'd23701; ROM4[9038]<=16'd57212;
ROM1[9039]<=16'd4789; ROM2[9039]<=16'd0; ROM3[9039]<=16'd23680; ROM4[9039]<=16'd57201;
ROM1[9040]<=16'd4803; ROM2[9040]<=16'd0; ROM3[9040]<=16'd23675; ROM4[9040]<=16'd57199;
ROM1[9041]<=16'd4814; ROM2[9041]<=16'd0; ROM3[9041]<=16'd23706; ROM4[9041]<=16'd57223;
ROM1[9042]<=16'd4814; ROM2[9042]<=16'd0; ROM3[9042]<=16'd23733; ROM4[9042]<=16'd57245;
ROM1[9043]<=16'd4786; ROM2[9043]<=16'd0; ROM3[9043]<=16'd23725; ROM4[9043]<=16'd57230;
ROM1[9044]<=16'd4755; ROM2[9044]<=16'd0; ROM3[9044]<=16'd23714; ROM4[9044]<=16'd57213;
ROM1[9045]<=16'd4743; ROM2[9045]<=16'd0; ROM3[9045]<=16'd23715; ROM4[9045]<=16'd57211;
ROM1[9046]<=16'd4749; ROM2[9046]<=16'd0; ROM3[9046]<=16'd23709; ROM4[9046]<=16'd57211;
ROM1[9047]<=16'd4787; ROM2[9047]<=16'd0; ROM3[9047]<=16'd23713; ROM4[9047]<=16'd57224;
ROM1[9048]<=16'd4818; ROM2[9048]<=16'd0; ROM3[9048]<=16'd23714; ROM4[9048]<=16'd57233;
ROM1[9049]<=16'd4814; ROM2[9049]<=16'd0; ROM3[9049]<=16'd23717; ROM4[9049]<=16'd57232;
ROM1[9050]<=16'd4797; ROM2[9050]<=16'd0; ROM3[9050]<=16'd23717; ROM4[9050]<=16'd57233;
ROM1[9051]<=16'd4781; ROM2[9051]<=16'd0; ROM3[9051]<=16'd23718; ROM4[9051]<=16'd57237;
ROM1[9052]<=16'd4769; ROM2[9052]<=16'd0; ROM3[9052]<=16'd23720; ROM4[9052]<=16'd57236;
ROM1[9053]<=16'd4771; ROM2[9053]<=16'd0; ROM3[9053]<=16'd23733; ROM4[9053]<=16'd57248;
ROM1[9054]<=16'd4788; ROM2[9054]<=16'd0; ROM3[9054]<=16'd23737; ROM4[9054]<=16'd57261;
ROM1[9055]<=16'd4789; ROM2[9055]<=16'd0; ROM3[9055]<=16'd23702; ROM4[9055]<=16'd57238;
ROM1[9056]<=16'd4804; ROM2[9056]<=16'd0; ROM3[9056]<=16'd23674; ROM4[9056]<=16'd57225;
ROM1[9057]<=16'd4816; ROM2[9057]<=16'd0; ROM3[9057]<=16'd23674; ROM4[9057]<=16'd57235;
ROM1[9058]<=16'd4801; ROM2[9058]<=16'd0; ROM3[9058]<=16'd23680; ROM4[9058]<=16'd57233;
ROM1[9059]<=16'd4789; ROM2[9059]<=16'd0; ROM3[9059]<=16'd23690; ROM4[9059]<=16'd57233;
ROM1[9060]<=16'd4779; ROM2[9060]<=16'd0; ROM3[9060]<=16'd23694; ROM4[9060]<=16'd57236;
ROM1[9061]<=16'd4757; ROM2[9061]<=16'd0; ROM3[9061]<=16'd23693; ROM4[9061]<=16'd57228;
ROM1[9062]<=16'd4753; ROM2[9062]<=16'd0; ROM3[9062]<=16'd23691; ROM4[9062]<=16'd57224;
ROM1[9063]<=16'd4788; ROM2[9063]<=16'd0; ROM3[9063]<=16'd23703; ROM4[9063]<=16'd57242;
ROM1[9064]<=16'd4822; ROM2[9064]<=16'd0; ROM3[9064]<=16'd23698; ROM4[9064]<=16'd57246;
ROM1[9065]<=16'd4819; ROM2[9065]<=16'd0; ROM3[9065]<=16'd23674; ROM4[9065]<=16'd57229;
ROM1[9066]<=16'd4804; ROM2[9066]<=16'd0; ROM3[9066]<=16'd23679; ROM4[9066]<=16'd57227;
ROM1[9067]<=16'd4804; ROM2[9067]<=16'd0; ROM3[9067]<=16'd23713; ROM4[9067]<=16'd57245;
ROM1[9068]<=16'd4789; ROM2[9068]<=16'd0; ROM3[9068]<=16'd23723; ROM4[9068]<=16'd57245;
ROM1[9069]<=16'd4759; ROM2[9069]<=16'd0; ROM3[9069]<=16'd23716; ROM4[9069]<=16'd57224;
ROM1[9070]<=16'd4752; ROM2[9070]<=16'd0; ROM3[9070]<=16'd23721; ROM4[9070]<=16'd57225;
ROM1[9071]<=16'd4754; ROM2[9071]<=16'd0; ROM3[9071]<=16'd23711; ROM4[9071]<=16'd57219;
ROM1[9072]<=16'd4787; ROM2[9072]<=16'd0; ROM3[9072]<=16'd23710; ROM4[9072]<=16'd57223;
ROM1[9073]<=16'd4824; ROM2[9073]<=16'd0; ROM3[9073]<=16'd23721; ROM4[9073]<=16'd57241;
ROM1[9074]<=16'd4809; ROM2[9074]<=16'd0; ROM3[9074]<=16'd23716; ROM4[9074]<=16'd57232;
ROM1[9075]<=16'd4786; ROM2[9075]<=16'd0; ROM3[9075]<=16'd23714; ROM4[9075]<=16'd57223;
ROM1[9076]<=16'd4778; ROM2[9076]<=16'd0; ROM3[9076]<=16'd23730; ROM4[9076]<=16'd57230;
ROM1[9077]<=16'd4769; ROM2[9077]<=16'd0; ROM3[9077]<=16'd23740; ROM4[9077]<=16'd57235;
ROM1[9078]<=16'd4753; ROM2[9078]<=16'd0; ROM3[9078]<=16'd23747; ROM4[9078]<=16'd57237;
ROM1[9079]<=16'd4759; ROM2[9079]<=16'd0; ROM3[9079]<=16'd23750; ROM4[9079]<=16'd57243;
ROM1[9080]<=16'd4791; ROM2[9080]<=16'd0; ROM3[9080]<=16'd23744; ROM4[9080]<=16'd57246;
ROM1[9081]<=16'd4832; ROM2[9081]<=16'd0; ROM3[9081]<=16'd23741; ROM4[9081]<=16'd57253;
ROM1[9082]<=16'd4844; ROM2[9082]<=16'd0; ROM3[9082]<=16'd23744; ROM4[9082]<=16'd57259;
ROM1[9083]<=16'd4825; ROM2[9083]<=16'd0; ROM3[9083]<=16'd23746; ROM4[9083]<=16'd57259;
ROM1[9084]<=16'd4803; ROM2[9084]<=16'd0; ROM3[9084]<=16'd23747; ROM4[9084]<=16'd57261;
ROM1[9085]<=16'd4795; ROM2[9085]<=16'd0; ROM3[9085]<=16'd23753; ROM4[9085]<=16'd57266;
ROM1[9086]<=16'd4785; ROM2[9086]<=16'd0; ROM3[9086]<=16'd23754; ROM4[9086]<=16'd57266;
ROM1[9087]<=16'd4788; ROM2[9087]<=16'd0; ROM3[9087]<=16'd23751; ROM4[9087]<=16'd57266;
ROM1[9088]<=16'd4807; ROM2[9088]<=16'd0; ROM3[9088]<=16'd23745; ROM4[9088]<=16'd57266;
ROM1[9089]<=16'd4833; ROM2[9089]<=16'd0; ROM3[9089]<=16'd23719; ROM4[9089]<=16'd57258;
ROM1[9090]<=16'd4838; ROM2[9090]<=16'd0; ROM3[9090]<=16'd23696; ROM4[9090]<=16'd57243;
ROM1[9091]<=16'd4833; ROM2[9091]<=16'd0; ROM3[9091]<=16'd23703; ROM4[9091]<=16'd57244;
ROM1[9092]<=16'd4841; ROM2[9092]<=16'd0; ROM3[9092]<=16'd23738; ROM4[9092]<=16'd57272;
ROM1[9093]<=16'd4821; ROM2[9093]<=16'd0; ROM3[9093]<=16'd23741; ROM4[9093]<=16'd57269;
ROM1[9094]<=16'd4780; ROM2[9094]<=16'd0; ROM3[9094]<=16'd23722; ROM4[9094]<=16'd57244;
ROM1[9095]<=16'd4788; ROM2[9095]<=16'd0; ROM3[9095]<=16'd23742; ROM4[9095]<=16'd57260;
ROM1[9096]<=16'd4798; ROM2[9096]<=16'd0; ROM3[9096]<=16'd23733; ROM4[9096]<=16'd57260;
ROM1[9097]<=16'd4801; ROM2[9097]<=16'd0; ROM3[9097]<=16'd23702; ROM4[9097]<=16'd57238;
ROM1[9098]<=16'd4820; ROM2[9098]<=16'd0; ROM3[9098]<=16'd23689; ROM4[9098]<=16'd57236;
ROM1[9099]<=16'd4803; ROM2[9099]<=16'd0; ROM3[9099]<=16'd23672; ROM4[9099]<=16'd57226;
ROM1[9100]<=16'd4774; ROM2[9100]<=16'd0; ROM3[9100]<=16'd23672; ROM4[9100]<=16'd57214;
ROM1[9101]<=16'd4770; ROM2[9101]<=16'd0; ROM3[9101]<=16'd23695; ROM4[9101]<=16'd57228;
ROM1[9102]<=16'd4773; ROM2[9102]<=16'd0; ROM3[9102]<=16'd23716; ROM4[9102]<=16'd57246;
ROM1[9103]<=16'd4758; ROM2[9103]<=16'd0; ROM3[9103]<=16'd23720; ROM4[9103]<=16'd57250;
ROM1[9104]<=16'd4766; ROM2[9104]<=16'd0; ROM3[9104]<=16'd23723; ROM4[9104]<=16'd57258;
ROM1[9105]<=16'd4791; ROM2[9105]<=16'd0; ROM3[9105]<=16'd23714; ROM4[9105]<=16'd57257;
ROM1[9106]<=16'd4805; ROM2[9106]<=16'd0; ROM3[9106]<=16'd23686; ROM4[9106]<=16'd57236;
ROM1[9107]<=16'd4800; ROM2[9107]<=16'd0; ROM3[9107]<=16'd23672; ROM4[9107]<=16'd57222;
ROM1[9108]<=16'd4778; ROM2[9108]<=16'd0; ROM3[9108]<=16'd23668; ROM4[9108]<=16'd57216;
ROM1[9109]<=16'd4766; ROM2[9109]<=16'd0; ROM3[9109]<=16'd23680; ROM4[9109]<=16'd57219;
ROM1[9110]<=16'd4764; ROM2[9110]<=16'd0; ROM3[9110]<=16'd23702; ROM4[9110]<=16'd57227;
ROM1[9111]<=16'd4750; ROM2[9111]<=16'd0; ROM3[9111]<=16'd23711; ROM4[9111]<=16'd57227;
ROM1[9112]<=16'd4746; ROM2[9112]<=16'd0; ROM3[9112]<=16'd23708; ROM4[9112]<=16'd57223;
ROM1[9113]<=16'd4765; ROM2[9113]<=16'd0; ROM3[9113]<=16'd23706; ROM4[9113]<=16'd57224;
ROM1[9114]<=16'd4803; ROM2[9114]<=16'd0; ROM3[9114]<=16'd23707; ROM4[9114]<=16'd57232;
ROM1[9115]<=16'd4816; ROM2[9115]<=16'd0; ROM3[9115]<=16'd23701; ROM4[9115]<=16'd57231;
ROM1[9116]<=16'd4799; ROM2[9116]<=16'd0; ROM3[9116]<=16'd23698; ROM4[9116]<=16'd57217;
ROM1[9117]<=16'd4779; ROM2[9117]<=16'd0; ROM3[9117]<=16'd23701; ROM4[9117]<=16'd57215;
ROM1[9118]<=16'd4773; ROM2[9118]<=16'd0; ROM3[9118]<=16'd23707; ROM4[9118]<=16'd57222;
ROM1[9119]<=16'd4760; ROM2[9119]<=16'd0; ROM3[9119]<=16'd23713; ROM4[9119]<=16'd57225;
ROM1[9120]<=16'd4751; ROM2[9120]<=16'd0; ROM3[9120]<=16'd23717; ROM4[9120]<=16'd57229;
ROM1[9121]<=16'd4762; ROM2[9121]<=16'd0; ROM3[9121]<=16'd23721; ROM4[9121]<=16'd57234;
ROM1[9122]<=16'd4791; ROM2[9122]<=16'd0; ROM3[9122]<=16'd23710; ROM4[9122]<=16'd57232;
ROM1[9123]<=16'd4810; ROM2[9123]<=16'd0; ROM3[9123]<=16'd23691; ROM4[9123]<=16'd57222;
ROM1[9124]<=16'd4796; ROM2[9124]<=16'd0; ROM3[9124]<=16'd23686; ROM4[9124]<=16'd57211;
ROM1[9125]<=16'd4790; ROM2[9125]<=16'd0; ROM3[9125]<=16'd23697; ROM4[9125]<=16'd57221;
ROM1[9126]<=16'd4790; ROM2[9126]<=16'd0; ROM3[9126]<=16'd23711; ROM4[9126]<=16'd57230;
ROM1[9127]<=16'd4776; ROM2[9127]<=16'd0; ROM3[9127]<=16'd23713; ROM4[9127]<=16'd57228;
ROM1[9128]<=16'd4760; ROM2[9128]<=16'd0; ROM3[9128]<=16'd23713; ROM4[9128]<=16'd57222;
ROM1[9129]<=16'd4769; ROM2[9129]<=16'd0; ROM3[9129]<=16'd23715; ROM4[9129]<=16'd57222;
ROM1[9130]<=16'd4777; ROM2[9130]<=16'd0; ROM3[9130]<=16'd23696; ROM4[9130]<=16'd57212;
ROM1[9131]<=16'd4788; ROM2[9131]<=16'd0; ROM3[9131]<=16'd23664; ROM4[9131]<=16'd57191;
ROM1[9132]<=16'd4798; ROM2[9132]<=16'd0; ROM3[9132]<=16'd23661; ROM4[9132]<=16'd57194;
ROM1[9133]<=16'd4787; ROM2[9133]<=16'd0; ROM3[9133]<=16'd23668; ROM4[9133]<=16'd57201;
ROM1[9134]<=16'd4771; ROM2[9134]<=16'd0; ROM3[9134]<=16'd23683; ROM4[9134]<=16'd57208;
ROM1[9135]<=16'd4776; ROM2[9135]<=16'd0; ROM3[9135]<=16'd23702; ROM4[9135]<=16'd57224;
ROM1[9136]<=16'd4789; ROM2[9136]<=16'd0; ROM3[9136]<=16'd23729; ROM4[9136]<=16'd57249;
ROM1[9137]<=16'd4792; ROM2[9137]<=16'd0; ROM3[9137]<=16'd23736; ROM4[9137]<=16'd57254;
ROM1[9138]<=16'd4794; ROM2[9138]<=16'd0; ROM3[9138]<=16'd23721; ROM4[9138]<=16'd57241;
ROM1[9139]<=16'd4815; ROM2[9139]<=16'd0; ROM3[9139]<=16'd23701; ROM4[9139]<=16'd57237;
ROM1[9140]<=16'd4818; ROM2[9140]<=16'd0; ROM3[9140]<=16'd23682; ROM4[9140]<=16'd57228;
ROM1[9141]<=16'd4809; ROM2[9141]<=16'd0; ROM3[9141]<=16'd23684; ROM4[9141]<=16'd57224;
ROM1[9142]<=16'd4807; ROM2[9142]<=16'd0; ROM3[9142]<=16'd23707; ROM4[9142]<=16'd57239;
ROM1[9143]<=16'd4803; ROM2[9143]<=16'd0; ROM3[9143]<=16'd23731; ROM4[9143]<=16'd57252;
ROM1[9144]<=16'd4793; ROM2[9144]<=16'd0; ROM3[9144]<=16'd23742; ROM4[9144]<=16'd57258;
ROM1[9145]<=16'd4788; ROM2[9145]<=16'd0; ROM3[9145]<=16'd23746; ROM4[9145]<=16'd57260;
ROM1[9146]<=16'd4798; ROM2[9146]<=16'd0; ROM3[9146]<=16'd23743; ROM4[9146]<=16'd57258;
ROM1[9147]<=16'd4825; ROM2[9147]<=16'd0; ROM3[9147]<=16'd23735; ROM4[9147]<=16'd57255;
ROM1[9148]<=16'd4850; ROM2[9148]<=16'd0; ROM3[9148]<=16'd23732; ROM4[9148]<=16'd57259;
ROM1[9149]<=16'd4824; ROM2[9149]<=16'd0; ROM3[9149]<=16'd23711; ROM4[9149]<=16'd57241;
ROM1[9150]<=16'd4794; ROM2[9150]<=16'd0; ROM3[9150]<=16'd23703; ROM4[9150]<=16'd57230;
ROM1[9151]<=16'd4778; ROM2[9151]<=16'd0; ROM3[9151]<=16'd23711; ROM4[9151]<=16'd57230;
ROM1[9152]<=16'd4757; ROM2[9152]<=16'd0; ROM3[9152]<=16'd23707; ROM4[9152]<=16'd57224;
ROM1[9153]<=16'd4755; ROM2[9153]<=16'd0; ROM3[9153]<=16'd23722; ROM4[9153]<=16'd57234;
ROM1[9154]<=16'd4772; ROM2[9154]<=16'd0; ROM3[9154]<=16'd23729; ROM4[9154]<=16'd57243;
ROM1[9155]<=16'd4796; ROM2[9155]<=16'd0; ROM3[9155]<=16'd23713; ROM4[9155]<=16'd57237;
ROM1[9156]<=16'd4819; ROM2[9156]<=16'd0; ROM3[9156]<=16'd23695; ROM4[9156]<=16'd57230;
ROM1[9157]<=16'd4818; ROM2[9157]<=16'd0; ROM3[9157]<=16'd23686; ROM4[9157]<=16'd57226;
ROM1[9158]<=16'd4805; ROM2[9158]<=16'd0; ROM3[9158]<=16'd23692; ROM4[9158]<=16'd57230;
ROM1[9159]<=16'd4792; ROM2[9159]<=16'd0; ROM3[9159]<=16'd23704; ROM4[9159]<=16'd57232;
ROM1[9160]<=16'd4780; ROM2[9160]<=16'd0; ROM3[9160]<=16'd23711; ROM4[9160]<=16'd57233;
ROM1[9161]<=16'd4772; ROM2[9161]<=16'd0; ROM3[9161]<=16'd23722; ROM4[9161]<=16'd57237;
ROM1[9162]<=16'd4778; ROM2[9162]<=16'd0; ROM3[9162]<=16'd23727; ROM4[9162]<=16'd57241;
ROM1[9163]<=16'd4795; ROM2[9163]<=16'd0; ROM3[9163]<=16'd23718; ROM4[9163]<=16'd57238;
ROM1[9164]<=16'd4813; ROM2[9164]<=16'd0; ROM3[9164]<=16'd23698; ROM4[9164]<=16'd57224;
ROM1[9165]<=16'd4818; ROM2[9165]<=16'd0; ROM3[9165]<=16'd23683; ROM4[9165]<=16'd57216;
ROM1[9166]<=16'd4805; ROM2[9166]<=16'd0; ROM3[9166]<=16'd23684; ROM4[9166]<=16'd57210;
ROM1[9167]<=16'd4781; ROM2[9167]<=16'd0; ROM3[9167]<=16'd23692; ROM4[9167]<=16'd57210;
ROM1[9168]<=16'd4769; ROM2[9168]<=16'd0; ROM3[9168]<=16'd23697; ROM4[9168]<=16'd57210;
ROM1[9169]<=16'd4753; ROM2[9169]<=16'd0; ROM3[9169]<=16'd23700; ROM4[9169]<=16'd57204;
ROM1[9170]<=16'd4761; ROM2[9170]<=16'd0; ROM3[9170]<=16'd23720; ROM4[9170]<=16'd57225;
ROM1[9171]<=16'd4789; ROM2[9171]<=16'd0; ROM3[9171]<=16'd23727; ROM4[9171]<=16'd57243;
ROM1[9172]<=16'd4798; ROM2[9172]<=16'd0; ROM3[9172]<=16'd23703; ROM4[9172]<=16'd57225;
ROM1[9173]<=16'd4804; ROM2[9173]<=16'd0; ROM3[9173]<=16'd23679; ROM4[9173]<=16'd57213;
ROM1[9174]<=16'd4784; ROM2[9174]<=16'd0; ROM3[9174]<=16'd23664; ROM4[9174]<=16'd57198;
ROM1[9175]<=16'd4760; ROM2[9175]<=16'd0; ROM3[9175]<=16'd23665; ROM4[9175]<=16'd57189;
ROM1[9176]<=16'd4758; ROM2[9176]<=16'd0; ROM3[9176]<=16'd23680; ROM4[9176]<=16'd57199;
ROM1[9177]<=16'd4750; ROM2[9177]<=16'd0; ROM3[9177]<=16'd23689; ROM4[9177]<=16'd57200;
ROM1[9178]<=16'd4737; ROM2[9178]<=16'd0; ROM3[9178]<=16'd23691; ROM4[9178]<=16'd57200;
ROM1[9179]<=16'd4760; ROM2[9179]<=16'd0; ROM3[9179]<=16'd23707; ROM4[9179]<=16'd57217;
ROM1[9180]<=16'd4791; ROM2[9180]<=16'd0; ROM3[9180]<=16'd23704; ROM4[9180]<=16'd57222;
ROM1[9181]<=16'd4817; ROM2[9181]<=16'd0; ROM3[9181]<=16'd23684; ROM4[9181]<=16'd57216;
ROM1[9182]<=16'd4832; ROM2[9182]<=16'd0; ROM3[9182]<=16'd23691; ROM4[9182]<=16'd57223;
ROM1[9183]<=16'd4793; ROM2[9183]<=16'd0; ROM3[9183]<=16'd23676; ROM4[9183]<=16'd57198;
ROM1[9184]<=16'd4761; ROM2[9184]<=16'd0; ROM3[9184]<=16'd23672; ROM4[9184]<=16'd57187;
ROM1[9185]<=16'd4760; ROM2[9185]<=16'd0; ROM3[9185]<=16'd23689; ROM4[9185]<=16'd57198;
ROM1[9186]<=16'd4731; ROM2[9186]<=16'd0; ROM3[9186]<=16'd23678; ROM4[9186]<=16'd57186;
ROM1[9187]<=16'd4730; ROM2[9187]<=16'd0; ROM3[9187]<=16'd23680; ROM4[9187]<=16'd57189;
ROM1[9188]<=16'd4760; ROM2[9188]<=16'd0; ROM3[9188]<=16'd23688; ROM4[9188]<=16'd57197;
ROM1[9189]<=16'd4790; ROM2[9189]<=16'd0; ROM3[9189]<=16'd23674; ROM4[9189]<=16'd57199;
ROM1[9190]<=16'd4801; ROM2[9190]<=16'd0; ROM3[9190]<=16'd23665; ROM4[9190]<=16'd57197;
ROM1[9191]<=16'd4790; ROM2[9191]<=16'd0; ROM3[9191]<=16'd23668; ROM4[9191]<=16'd57194;
ROM1[9192]<=16'd4782; ROM2[9192]<=16'd0; ROM3[9192]<=16'd23686; ROM4[9192]<=16'd57208;
ROM1[9193]<=16'd4777; ROM2[9193]<=16'd0; ROM3[9193]<=16'd23706; ROM4[9193]<=16'd57223;
ROM1[9194]<=16'd4761; ROM2[9194]<=16'd0; ROM3[9194]<=16'd23712; ROM4[9194]<=16'd57218;
ROM1[9195]<=16'd4756; ROM2[9195]<=16'd0; ROM3[9195]<=16'd23708; ROM4[9195]<=16'd57218;
ROM1[9196]<=16'd4763; ROM2[9196]<=16'd0; ROM3[9196]<=16'd23697; ROM4[9196]<=16'd57213;
ROM1[9197]<=16'd4786; ROM2[9197]<=16'd0; ROM3[9197]<=16'd23684; ROM4[9197]<=16'd57207;
ROM1[9198]<=16'd4807; ROM2[9198]<=16'd0; ROM3[9198]<=16'd23673; ROM4[9198]<=16'd57210;
ROM1[9199]<=16'd4805; ROM2[9199]<=16'd0; ROM3[9199]<=16'd23680; ROM4[9199]<=16'd57216;
ROM1[9200]<=16'd4796; ROM2[9200]<=16'd0; ROM3[9200]<=16'd23691; ROM4[9200]<=16'd57223;
ROM1[9201]<=16'd4787; ROM2[9201]<=16'd0; ROM3[9201]<=16'd23704; ROM4[9201]<=16'd57226;
ROM1[9202]<=16'd4782; ROM2[9202]<=16'd0; ROM3[9202]<=16'd23717; ROM4[9202]<=16'd57236;
ROM1[9203]<=16'd4773; ROM2[9203]<=16'd0; ROM3[9203]<=16'd23723; ROM4[9203]<=16'd57239;
ROM1[9204]<=16'd4776; ROM2[9204]<=16'd0; ROM3[9204]<=16'd23724; ROM4[9204]<=16'd57242;
ROM1[9205]<=16'd4801; ROM2[9205]<=16'd0; ROM3[9205]<=16'd23715; ROM4[9205]<=16'd57244;
ROM1[9206]<=16'd4833; ROM2[9206]<=16'd0; ROM3[9206]<=16'd23707; ROM4[9206]<=16'd57244;
ROM1[9207]<=16'd4841; ROM2[9207]<=16'd0; ROM3[9207]<=16'd23714; ROM4[9207]<=16'd57250;
ROM1[9208]<=16'd4822; ROM2[9208]<=16'd0; ROM3[9208]<=16'd23722; ROM4[9208]<=16'd57249;
ROM1[9209]<=16'd4815; ROM2[9209]<=16'd0; ROM3[9209]<=16'd23744; ROM4[9209]<=16'd57260;
ROM1[9210]<=16'd4810; ROM2[9210]<=16'd0; ROM3[9210]<=16'd23759; ROM4[9210]<=16'd57269;
ROM1[9211]<=16'd4775; ROM2[9211]<=16'd0; ROM3[9211]<=16'd23749; ROM4[9211]<=16'd57251;
ROM1[9212]<=16'd4767; ROM2[9212]<=16'd0; ROM3[9212]<=16'd23742; ROM4[9212]<=16'd57243;
ROM1[9213]<=16'd4790; ROM2[9213]<=16'd0; ROM3[9213]<=16'd23738; ROM4[9213]<=16'd57248;
ROM1[9214]<=16'd4820; ROM2[9214]<=16'd0; ROM3[9214]<=16'd23729; ROM4[9214]<=16'd57247;
ROM1[9215]<=16'd4834; ROM2[9215]<=16'd0; ROM3[9215]<=16'd23731; ROM4[9215]<=16'd57254;
ROM1[9216]<=16'd4821; ROM2[9216]<=16'd0; ROM3[9216]<=16'd23734; ROM4[9216]<=16'd57253;
ROM1[9217]<=16'd4800; ROM2[9217]<=16'd0; ROM3[9217]<=16'd23742; ROM4[9217]<=16'd57251;
ROM1[9218]<=16'd4782; ROM2[9218]<=16'd0; ROM3[9218]<=16'd23744; ROM4[9218]<=16'd57249;
ROM1[9219]<=16'd4769; ROM2[9219]<=16'd0; ROM3[9219]<=16'd23741; ROM4[9219]<=16'd57243;
ROM1[9220]<=16'd4767; ROM2[9220]<=16'd0; ROM3[9220]<=16'd23744; ROM4[9220]<=16'd57245;
ROM1[9221]<=16'd4770; ROM2[9221]<=16'd0; ROM3[9221]<=16'd23732; ROM4[9221]<=16'd57237;
ROM1[9222]<=16'd4793; ROM2[9222]<=16'd0; ROM3[9222]<=16'd23716; ROM4[9222]<=16'd57231;
ROM1[9223]<=16'd4822; ROM2[9223]<=16'd0; ROM3[9223]<=16'd23712; ROM4[9223]<=16'd57240;
ROM1[9224]<=16'd4826; ROM2[9224]<=16'd0; ROM3[9224]<=16'd23721; ROM4[9224]<=16'd57247;
ROM1[9225]<=16'd4798; ROM2[9225]<=16'd0; ROM3[9225]<=16'd23716; ROM4[9225]<=16'd57237;
ROM1[9226]<=16'd4763; ROM2[9226]<=16'd0; ROM3[9226]<=16'd23711; ROM4[9226]<=16'd57226;
ROM1[9227]<=16'd4747; ROM2[9227]<=16'd0; ROM3[9227]<=16'd23715; ROM4[9227]<=16'd57220;
ROM1[9228]<=16'd4733; ROM2[9228]<=16'd0; ROM3[9228]<=16'd23712; ROM4[9228]<=16'd57217;
ROM1[9229]<=16'd4743; ROM2[9229]<=16'd0; ROM3[9229]<=16'd23717; ROM4[9229]<=16'd57229;
ROM1[9230]<=16'd4781; ROM2[9230]<=16'd0; ROM3[9230]<=16'd23723; ROM4[9230]<=16'd57244;
ROM1[9231]<=16'd4808; ROM2[9231]<=16'd0; ROM3[9231]<=16'd23704; ROM4[9231]<=16'd57238;
ROM1[9232]<=16'd4812; ROM2[9232]<=16'd0; ROM3[9232]<=16'd23705; ROM4[9232]<=16'd57239;
ROM1[9233]<=16'd4799; ROM2[9233]<=16'd0; ROM3[9233]<=16'd23716; ROM4[9233]<=16'd57239;
ROM1[9234]<=16'd4770; ROM2[9234]<=16'd0; ROM3[9234]<=16'd23703; ROM4[9234]<=16'd57222;
ROM1[9235]<=16'd4767; ROM2[9235]<=16'd0; ROM3[9235]<=16'd23714; ROM4[9235]<=16'd57232;
ROM1[9236]<=16'd4746; ROM2[9236]<=16'd0; ROM3[9236]<=16'd23717; ROM4[9236]<=16'd57227;
ROM1[9237]<=16'd4733; ROM2[9237]<=16'd0; ROM3[9237]<=16'd23704; ROM4[9237]<=16'd57213;
ROM1[9238]<=16'd4755; ROM2[9238]<=16'd0; ROM3[9238]<=16'd23701; ROM4[9238]<=16'd57215;
ROM1[9239]<=16'd4780; ROM2[9239]<=16'd0; ROM3[9239]<=16'd23685; ROM4[9239]<=16'd57214;
ROM1[9240]<=16'd4786; ROM2[9240]<=16'd0; ROM3[9240]<=16'd23667; ROM4[9240]<=16'd57204;
ROM1[9241]<=16'd4766; ROM2[9241]<=16'd0; ROM3[9241]<=16'd23660; ROM4[9241]<=16'd57192;
ROM1[9242]<=16'd4749; ROM2[9242]<=16'd0; ROM3[9242]<=16'd23670; ROM4[9242]<=16'd57189;
ROM1[9243]<=16'd4747; ROM2[9243]<=16'd0; ROM3[9243]<=16'd23685; ROM4[9243]<=16'd57198;
ROM1[9244]<=16'd4740; ROM2[9244]<=16'd0; ROM3[9244]<=16'd23701; ROM4[9244]<=16'd57208;
ROM1[9245]<=16'd4741; ROM2[9245]<=16'd0; ROM3[9245]<=16'd23708; ROM4[9245]<=16'd57212;
ROM1[9246]<=16'd4754; ROM2[9246]<=16'd0; ROM3[9246]<=16'd23705; ROM4[9246]<=16'd57216;
ROM1[9247]<=16'd4784; ROM2[9247]<=16'd0; ROM3[9247]<=16'd23697; ROM4[9247]<=16'd57215;
ROM1[9248]<=16'd4821; ROM2[9248]<=16'd0; ROM3[9248]<=16'd23699; ROM4[9248]<=16'd57227;
ROM1[9249]<=16'd4806; ROM2[9249]<=16'd0; ROM3[9249]<=16'd23696; ROM4[9249]<=16'd57221;
ROM1[9250]<=16'd4777; ROM2[9250]<=16'd0; ROM3[9250]<=16'd23693; ROM4[9250]<=16'd57212;
ROM1[9251]<=16'd4761; ROM2[9251]<=16'd0; ROM3[9251]<=16'd23704; ROM4[9251]<=16'd57213;
ROM1[9252]<=16'd4747; ROM2[9252]<=16'd0; ROM3[9252]<=16'd23707; ROM4[9252]<=16'd57209;
ROM1[9253]<=16'd4749; ROM2[9253]<=16'd0; ROM3[9253]<=16'd23724; ROM4[9253]<=16'd57222;
ROM1[9254]<=16'd4761; ROM2[9254]<=16'd0; ROM3[9254]<=16'd23735; ROM4[9254]<=16'd57233;
ROM1[9255]<=16'd4776; ROM2[9255]<=16'd0; ROM3[9255]<=16'd23721; ROM4[9255]<=16'd57225;
ROM1[9256]<=16'd4798; ROM2[9256]<=16'd0; ROM3[9256]<=16'd23705; ROM4[9256]<=16'd57218;
ROM1[9257]<=16'd4805; ROM2[9257]<=16'd0; ROM3[9257]<=16'd23703; ROM4[9257]<=16'd57223;
ROM1[9258]<=16'd4803; ROM2[9258]<=16'd0; ROM3[9258]<=16'd23715; ROM4[9258]<=16'd57233;
ROM1[9259]<=16'd4800; ROM2[9259]<=16'd0; ROM3[9259]<=16'd23729; ROM4[9259]<=16'd57241;
ROM1[9260]<=16'd4785; ROM2[9260]<=16'd0; ROM3[9260]<=16'd23731; ROM4[9260]<=16'd57244;
ROM1[9261]<=16'd4762; ROM2[9261]<=16'd0; ROM3[9261]<=16'd23725; ROM4[9261]<=16'd57231;
ROM1[9262]<=16'd4765; ROM2[9262]<=16'd0; ROM3[9262]<=16'd23723; ROM4[9262]<=16'd57235;
ROM1[9263]<=16'd4786; ROM2[9263]<=16'd0; ROM3[9263]<=16'd23720; ROM4[9263]<=16'd57246;
ROM1[9264]<=16'd4824; ROM2[9264]<=16'd0; ROM3[9264]<=16'd23711; ROM4[9264]<=16'd57250;
ROM1[9265]<=16'd4848; ROM2[9265]<=16'd0; ROM3[9265]<=16'd23716; ROM4[9265]<=16'd57265;
ROM1[9266]<=16'd4819; ROM2[9266]<=16'd0; ROM3[9266]<=16'd23709; ROM4[9266]<=16'd57254;
ROM1[9267]<=16'd4788; ROM2[9267]<=16'd0; ROM3[9267]<=16'd23704; ROM4[9267]<=16'd57242;
ROM1[9268]<=16'd4780; ROM2[9268]<=16'd0; ROM3[9268]<=16'd23720; ROM4[9268]<=16'd57252;
ROM1[9269]<=16'd4772; ROM2[9269]<=16'd0; ROM3[9269]<=16'd23731; ROM4[9269]<=16'd57255;
ROM1[9270]<=16'd4765; ROM2[9270]<=16'd0; ROM3[9270]<=16'd23730; ROM4[9270]<=16'd57250;
ROM1[9271]<=16'd4767; ROM2[9271]<=16'd0; ROM3[9271]<=16'd23720; ROM4[9271]<=16'd57241;
ROM1[9272]<=16'd4784; ROM2[9272]<=16'd0; ROM3[9272]<=16'd23703; ROM4[9272]<=16'd57227;
ROM1[9273]<=16'd4803; ROM2[9273]<=16'd0; ROM3[9273]<=16'd23689; ROM4[9273]<=16'd57222;
ROM1[9274]<=16'd4810; ROM2[9274]<=16'd0; ROM3[9274]<=16'd23702; ROM4[9274]<=16'd57230;
ROM1[9275]<=16'd4804; ROM2[9275]<=16'd0; ROM3[9275]<=16'd23723; ROM4[9275]<=16'd57238;
ROM1[9276]<=16'd4787; ROM2[9276]<=16'd0; ROM3[9276]<=16'd23730; ROM4[9276]<=16'd57239;
ROM1[9277]<=16'd4764; ROM2[9277]<=16'd0; ROM3[9277]<=16'd23726; ROM4[9277]<=16'd57232;
ROM1[9278]<=16'd4748; ROM2[9278]<=16'd0; ROM3[9278]<=16'd23729; ROM4[9278]<=16'd57229;
ROM1[9279]<=16'd4748; ROM2[9279]<=16'd0; ROM3[9279]<=16'd23720; ROM4[9279]<=16'd57222;
ROM1[9280]<=16'd4763; ROM2[9280]<=16'd0; ROM3[9280]<=16'd23703; ROM4[9280]<=16'd57212;
ROM1[9281]<=16'd4788; ROM2[9281]<=16'd0; ROM3[9281]<=16'd23690; ROM4[9281]<=16'd57209;
ROM1[9282]<=16'd4786; ROM2[9282]<=16'd0; ROM3[9282]<=16'd23683; ROM4[9282]<=16'd57203;
ROM1[9283]<=16'd4777; ROM2[9283]<=16'd0; ROM3[9283]<=16'd23694; ROM4[9283]<=16'd57209;
ROM1[9284]<=16'd4759; ROM2[9284]<=16'd0; ROM3[9284]<=16'd23705; ROM4[9284]<=16'd57213;
ROM1[9285]<=16'd4749; ROM2[9285]<=16'd0; ROM3[9285]<=16'd23719; ROM4[9285]<=16'd57217;
ROM1[9286]<=16'd4737; ROM2[9286]<=16'd0; ROM3[9286]<=16'd23728; ROM4[9286]<=16'd57225;
ROM1[9287]<=16'd4730; ROM2[9287]<=16'd0; ROM3[9287]<=16'd23729; ROM4[9287]<=16'd57227;
ROM1[9288]<=16'd4761; ROM2[9288]<=16'd0; ROM3[9288]<=16'd23728; ROM4[9288]<=16'd57233;
ROM1[9289]<=16'd4798; ROM2[9289]<=16'd0; ROM3[9289]<=16'd23711; ROM4[9289]<=16'd57232;
ROM1[9290]<=16'd4814; ROM2[9290]<=16'd0; ROM3[9290]<=16'd23704; ROM4[9290]<=16'd57227;
ROM1[9291]<=16'd4819; ROM2[9291]<=16'd0; ROM3[9291]<=16'd23718; ROM4[9291]<=16'd57237;
ROM1[9292]<=16'd4806; ROM2[9292]<=16'd0; ROM3[9292]<=16'd23724; ROM4[9292]<=16'd57240;
ROM1[9293]<=16'd4787; ROM2[9293]<=16'd0; ROM3[9293]<=16'd23725; ROM4[9293]<=16'd57237;
ROM1[9294]<=16'd4758; ROM2[9294]<=16'd0; ROM3[9294]<=16'd23711; ROM4[9294]<=16'd57219;
ROM1[9295]<=16'd4731; ROM2[9295]<=16'd0; ROM3[9295]<=16'd23688; ROM4[9295]<=16'd57193;
ROM1[9296]<=16'd4738; ROM2[9296]<=16'd0; ROM3[9296]<=16'd23673; ROM4[9296]<=16'd57180;
ROM1[9297]<=16'd4777; ROM2[9297]<=16'd0; ROM3[9297]<=16'd23667; ROM4[9297]<=16'd57186;
ROM1[9298]<=16'd4804; ROM2[9298]<=16'd0; ROM3[9298]<=16'd23664; ROM4[9298]<=16'd57192;
ROM1[9299]<=16'd4808; ROM2[9299]<=16'd0; ROM3[9299]<=16'd23673; ROM4[9299]<=16'd57204;
ROM1[9300]<=16'd4806; ROM2[9300]<=16'd0; ROM3[9300]<=16'd23693; ROM4[9300]<=16'd57222;
ROM1[9301]<=16'd4774; ROM2[9301]<=16'd0; ROM3[9301]<=16'd23684; ROM4[9301]<=16'd57209;
ROM1[9302]<=16'd4758; ROM2[9302]<=16'd0; ROM3[9302]<=16'd23686; ROM4[9302]<=16'd57207;
ROM1[9303]<=16'd4759; ROM2[9303]<=16'd0; ROM3[9303]<=16'd23704; ROM4[9303]<=16'd57217;
ROM1[9304]<=16'd4751; ROM2[9304]<=16'd0; ROM3[9304]<=16'd23690; ROM4[9304]<=16'd57204;
ROM1[9305]<=16'd4773; ROM2[9305]<=16'd0; ROM3[9305]<=16'd23681; ROM4[9305]<=16'd57204;
ROM1[9306]<=16'd4816; ROM2[9306]<=16'd0; ROM3[9306]<=16'd23685; ROM4[9306]<=16'd57218;
ROM1[9307]<=16'd4837; ROM2[9307]<=16'd0; ROM3[9307]<=16'd23697; ROM4[9307]<=16'd57236;
ROM1[9308]<=16'd4813; ROM2[9308]<=16'd0; ROM3[9308]<=16'd23697; ROM4[9308]<=16'd57228;
ROM1[9309]<=16'd4782; ROM2[9309]<=16'd0; ROM3[9309]<=16'd23691; ROM4[9309]<=16'd57217;
ROM1[9310]<=16'd4781; ROM2[9310]<=16'd0; ROM3[9310]<=16'd23706; ROM4[9310]<=16'd57227;
ROM1[9311]<=16'd4759; ROM2[9311]<=16'd0; ROM3[9311]<=16'd23706; ROM4[9311]<=16'd57217;
ROM1[9312]<=16'd4751; ROM2[9312]<=16'd0; ROM3[9312]<=16'd23698; ROM4[9312]<=16'd57211;
ROM1[9313]<=16'd4785; ROM2[9313]<=16'd0; ROM3[9313]<=16'd23709; ROM4[9313]<=16'd57225;
ROM1[9314]<=16'd4810; ROM2[9314]<=16'd0; ROM3[9314]<=16'd23697; ROM4[9314]<=16'd57218;
ROM1[9315]<=16'd4804; ROM2[9315]<=16'd0; ROM3[9315]<=16'd23672; ROM4[9315]<=16'd57203;
ROM1[9316]<=16'd4791; ROM2[9316]<=16'd0; ROM3[9316]<=16'd23675; ROM4[9316]<=16'd57202;
ROM1[9317]<=16'd4779; ROM2[9317]<=16'd0; ROM3[9317]<=16'd23696; ROM4[9317]<=16'd57210;
ROM1[9318]<=16'd4766; ROM2[9318]<=16'd0; ROM3[9318]<=16'd23697; ROM4[9318]<=16'd57209;
ROM1[9319]<=16'd4749; ROM2[9319]<=16'd0; ROM3[9319]<=16'd23698; ROM4[9319]<=16'd57204;
ROM1[9320]<=16'd4744; ROM2[9320]<=16'd0; ROM3[9320]<=16'd23708; ROM4[9320]<=16'd57212;
ROM1[9321]<=16'd4760; ROM2[9321]<=16'd0; ROM3[9321]<=16'd23711; ROM4[9321]<=16'd57220;
ROM1[9322]<=16'd4794; ROM2[9322]<=16'd0; ROM3[9322]<=16'd23711; ROM4[9322]<=16'd57226;
ROM1[9323]<=16'd4803; ROM2[9323]<=16'd0; ROM3[9323]<=16'd23694; ROM4[9323]<=16'd57217;
ROM1[9324]<=16'd4788; ROM2[9324]<=16'd0; ROM3[9324]<=16'd23685; ROM4[9324]<=16'd57207;
ROM1[9325]<=16'd4773; ROM2[9325]<=16'd0; ROM3[9325]<=16'd23696; ROM4[9325]<=16'd57212;
ROM1[9326]<=16'd4753; ROM2[9326]<=16'd0; ROM3[9326]<=16'd23699; ROM4[9326]<=16'd57208;
ROM1[9327]<=16'd4742; ROM2[9327]<=16'd0; ROM3[9327]<=16'd23705; ROM4[9327]<=16'd57208;
ROM1[9328]<=16'd4739; ROM2[9328]<=16'd0; ROM3[9328]<=16'd23714; ROM4[9328]<=16'd57218;
ROM1[9329]<=16'd4747; ROM2[9329]<=16'd0; ROM3[9329]<=16'd23713; ROM4[9329]<=16'd57219;
ROM1[9330]<=16'd4771; ROM2[9330]<=16'd0; ROM3[9330]<=16'd23702; ROM4[9330]<=16'd57218;
ROM1[9331]<=16'd4804; ROM2[9331]<=16'd0; ROM3[9331]<=16'd23696; ROM4[9331]<=16'd57222;
ROM1[9332]<=16'd4819; ROM2[9332]<=16'd0; ROM3[9332]<=16'd23708; ROM4[9332]<=16'd57232;
ROM1[9333]<=16'd4809; ROM2[9333]<=16'd0; ROM3[9333]<=16'd23719; ROM4[9333]<=16'd57237;
ROM1[9334]<=16'd4777; ROM2[9334]<=16'd0; ROM3[9334]<=16'd23711; ROM4[9334]<=16'd57222;
ROM1[9335]<=16'd4769; ROM2[9335]<=16'd0; ROM3[9335]<=16'd23719; ROM4[9335]<=16'd57229;
ROM1[9336]<=16'd4758; ROM2[9336]<=16'd0; ROM3[9336]<=16'd23729; ROM4[9336]<=16'd57235;
ROM1[9337]<=16'd4756; ROM2[9337]<=16'd0; ROM3[9337]<=16'd23725; ROM4[9337]<=16'd57232;
ROM1[9338]<=16'd4794; ROM2[9338]<=16'd0; ROM3[9338]<=16'd23740; ROM4[9338]<=16'd57252;
ROM1[9339]<=16'd4838; ROM2[9339]<=16'd0; ROM3[9339]<=16'd23746; ROM4[9339]<=16'd57265;
ROM1[9340]<=16'd4837; ROM2[9340]<=16'd0; ROM3[9340]<=16'd23723; ROM4[9340]<=16'd57250;
ROM1[9341]<=16'd4803; ROM2[9341]<=16'd0; ROM3[9341]<=16'd23704; ROM4[9341]<=16'd57224;
ROM1[9342]<=16'd4784; ROM2[9342]<=16'd0; ROM3[9342]<=16'd23710; ROM4[9342]<=16'd57221;
ROM1[9343]<=16'd4779; ROM2[9343]<=16'd0; ROM3[9343]<=16'd23724; ROM4[9343]<=16'd57232;
ROM1[9344]<=16'd4783; ROM2[9344]<=16'd0; ROM3[9344]<=16'd23745; ROM4[9344]<=16'd57245;
ROM1[9345]<=16'd4772; ROM2[9345]<=16'd0; ROM3[9345]<=16'd23743; ROM4[9345]<=16'd57241;
ROM1[9346]<=16'd4767; ROM2[9346]<=16'd0; ROM3[9346]<=16'd23724; ROM4[9346]<=16'd57226;
ROM1[9347]<=16'd4787; ROM2[9347]<=16'd0; ROM3[9347]<=16'd23705; ROM4[9347]<=16'd57214;
ROM1[9348]<=16'd4815; ROM2[9348]<=16'd0; ROM3[9348]<=16'd23700; ROM4[9348]<=16'd57223;
ROM1[9349]<=16'd4826; ROM2[9349]<=16'd0; ROM3[9349]<=16'd23718; ROM4[9349]<=16'd57242;
ROM1[9350]<=16'd4821; ROM2[9350]<=16'd0; ROM3[9350]<=16'd23734; ROM4[9350]<=16'd57253;
ROM1[9351]<=16'd4803; ROM2[9351]<=16'd0; ROM3[9351]<=16'd23742; ROM4[9351]<=16'd57254;
ROM1[9352]<=16'd4786; ROM2[9352]<=16'd0; ROM3[9352]<=16'd23746; ROM4[9352]<=16'd57252;
ROM1[9353]<=16'd4764; ROM2[9353]<=16'd0; ROM3[9353]<=16'd23738; ROM4[9353]<=16'd57243;
ROM1[9354]<=16'd4761; ROM2[9354]<=16'd0; ROM3[9354]<=16'd23727; ROM4[9354]<=16'd57235;
ROM1[9355]<=16'd4780; ROM2[9355]<=16'd0; ROM3[9355]<=16'd23711; ROM4[9355]<=16'd57227;
ROM1[9356]<=16'd4805; ROM2[9356]<=16'd0; ROM3[9356]<=16'd23695; ROM4[9356]<=16'd57220;
ROM1[9357]<=16'd4827; ROM2[9357]<=16'd0; ROM3[9357]<=16'd23712; ROM4[9357]<=16'd57238;
ROM1[9358]<=16'd4813; ROM2[9358]<=16'd0; ROM3[9358]<=16'd23723; ROM4[9358]<=16'd57249;
ROM1[9359]<=16'd4787; ROM2[9359]<=16'd0; ROM3[9359]<=16'd23724; ROM4[9359]<=16'd57243;
ROM1[9360]<=16'd4771; ROM2[9360]<=16'd0; ROM3[9360]<=16'd23728; ROM4[9360]<=16'd57244;
ROM1[9361]<=16'd4749; ROM2[9361]<=16'd0; ROM3[9361]<=16'd23723; ROM4[9361]<=16'd57232;
ROM1[9362]<=16'd4755; ROM2[9362]<=16'd0; ROM3[9362]<=16'd23726; ROM4[9362]<=16'd57235;
ROM1[9363]<=16'd4784; ROM2[9363]<=16'd0; ROM3[9363]<=16'd23724; ROM4[9363]<=16'd57242;
ROM1[9364]<=16'd4815; ROM2[9364]<=16'd0; ROM3[9364]<=16'd23708; ROM4[9364]<=16'd57234;
ROM1[9365]<=16'd4825; ROM2[9365]<=16'd0; ROM3[9365]<=16'd23695; ROM4[9365]<=16'd57230;
ROM1[9366]<=16'd4808; ROM2[9366]<=16'd0; ROM3[9366]<=16'd23690; ROM4[9366]<=16'd57221;
ROM1[9367]<=16'd4786; ROM2[9367]<=16'd0; ROM3[9367]<=16'd23691; ROM4[9367]<=16'd57212;
ROM1[9368]<=16'd4778; ROM2[9368]<=16'd0; ROM3[9368]<=16'd23697; ROM4[9368]<=16'd57216;
ROM1[9369]<=16'd4767; ROM2[9369]<=16'd0; ROM3[9369]<=16'd23707; ROM4[9369]<=16'd57216;
ROM1[9370]<=16'd4763; ROM2[9370]<=16'd0; ROM3[9370]<=16'd23710; ROM4[9370]<=16'd57217;
ROM1[9371]<=16'd4766; ROM2[9371]<=16'd0; ROM3[9371]<=16'd23697; ROM4[9371]<=16'd57210;
ROM1[9372]<=16'd4780; ROM2[9372]<=16'd0; ROM3[9372]<=16'd23670; ROM4[9372]<=16'd57195;
ROM1[9373]<=16'd4791; ROM2[9373]<=16'd0; ROM3[9373]<=16'd23650; ROM4[9373]<=16'd57188;
ROM1[9374]<=16'd4780; ROM2[9374]<=16'd0; ROM3[9374]<=16'd23650; ROM4[9374]<=16'd57187;
ROM1[9375]<=16'd4772; ROM2[9375]<=16'd0; ROM3[9375]<=16'd23663; ROM4[9375]<=16'd57195;
ROM1[9376]<=16'd4755; ROM2[9376]<=16'd0; ROM3[9376]<=16'd23670; ROM4[9376]<=16'd57197;
ROM1[9377]<=16'd4746; ROM2[9377]<=16'd0; ROM3[9377]<=16'd23687; ROM4[9377]<=16'd57206;
ROM1[9378]<=16'd4733; ROM2[9378]<=16'd0; ROM3[9378]<=16'd23694; ROM4[9378]<=16'd57206;
ROM1[9379]<=16'd4733; ROM2[9379]<=16'd0; ROM3[9379]<=16'd23694; ROM4[9379]<=16'd57201;
ROM1[9380]<=16'd4764; ROM2[9380]<=16'd0; ROM3[9380]<=16'd23697; ROM4[9380]<=16'd57210;
ROM1[9381]<=16'd4787; ROM2[9381]<=16'd0; ROM3[9381]<=16'd23679; ROM4[9381]<=16'd57205;
ROM1[9382]<=16'd4760; ROM2[9382]<=16'd0; ROM3[9382]<=16'd23651; ROM4[9382]<=16'd57178;
ROM1[9383]<=16'd4733; ROM2[9383]<=16'd0; ROM3[9383]<=16'd23652; ROM4[9383]<=16'd57167;
ROM1[9384]<=16'd4734; ROM2[9384]<=16'd0; ROM3[9384]<=16'd23687; ROM4[9384]<=16'd57185;
ROM1[9385]<=16'd4740; ROM2[9385]<=16'd0; ROM3[9385]<=16'd23714; ROM4[9385]<=16'd57203;
ROM1[9386]<=16'd4752; ROM2[9386]<=16'd0; ROM3[9386]<=16'd23742; ROM4[9386]<=16'd57228;
ROM1[9387]<=16'd4773; ROM2[9387]<=16'd0; ROM3[9387]<=16'd23758; ROM4[9387]<=16'd57246;
ROM1[9388]<=16'd4787; ROM2[9388]<=16'd0; ROM3[9388]<=16'd23747; ROM4[9388]<=16'd57239;
ROM1[9389]<=16'd4816; ROM2[9389]<=16'd0; ROM3[9389]<=16'd23734; ROM4[9389]<=16'd57236;
ROM1[9390]<=16'd4827; ROM2[9390]<=16'd0; ROM3[9390]<=16'd23727; ROM4[9390]<=16'd57232;
ROM1[9391]<=16'd4812; ROM2[9391]<=16'd0; ROM3[9391]<=16'd23729; ROM4[9391]<=16'd57232;
ROM1[9392]<=16'd4810; ROM2[9392]<=16'd0; ROM3[9392]<=16'd23748; ROM4[9392]<=16'd57250;
ROM1[9393]<=16'd4799; ROM2[9393]<=16'd0; ROM3[9393]<=16'd23750; ROM4[9393]<=16'd57246;
ROM1[9394]<=16'd4782; ROM2[9394]<=16'd0; ROM3[9394]<=16'd23746; ROM4[9394]<=16'd57240;
ROM1[9395]<=16'd4779; ROM2[9395]<=16'd0; ROM3[9395]<=16'd23749; ROM4[9395]<=16'd57244;
ROM1[9396]<=16'd4797; ROM2[9396]<=16'd0; ROM3[9396]<=16'd23748; ROM4[9396]<=16'd57255;
ROM1[9397]<=16'd4816; ROM2[9397]<=16'd0; ROM3[9397]<=16'd23724; ROM4[9397]<=16'd57247;
ROM1[9398]<=16'd4831; ROM2[9398]<=16'd0; ROM3[9398]<=16'd23704; ROM4[9398]<=16'd57237;
ROM1[9399]<=16'd4825; ROM2[9399]<=16'd0; ROM3[9399]<=16'd23702; ROM4[9399]<=16'd57237;
ROM1[9400]<=16'd4789; ROM2[9400]<=16'd0; ROM3[9400]<=16'd23692; ROM4[9400]<=16'd57214;
ROM1[9401]<=16'd4770; ROM2[9401]<=16'd0; ROM3[9401]<=16'd23700; ROM4[9401]<=16'd57209;
ROM1[9402]<=16'd4762; ROM2[9402]<=16'd0; ROM3[9402]<=16'd23716; ROM4[9402]<=16'd57219;
ROM1[9403]<=16'd4744; ROM2[9403]<=16'd0; ROM3[9403]<=16'd23712; ROM4[9403]<=16'd57212;
ROM1[9404]<=16'd4752; ROM2[9404]<=16'd0; ROM3[9404]<=16'd23714; ROM4[9404]<=16'd57211;
ROM1[9405]<=16'd4778; ROM2[9405]<=16'd0; ROM3[9405]<=16'd23710; ROM4[9405]<=16'd57216;
ROM1[9406]<=16'd4803; ROM2[9406]<=16'd0; ROM3[9406]<=16'd23695; ROM4[9406]<=16'd57214;
ROM1[9407]<=16'd4808; ROM2[9407]<=16'd0; ROM3[9407]<=16'd23701; ROM4[9407]<=16'd57221;
ROM1[9408]<=16'd4801; ROM2[9408]<=16'd0; ROM3[9408]<=16'd23716; ROM4[9408]<=16'd57230;
ROM1[9409]<=16'd4786; ROM2[9409]<=16'd0; ROM3[9409]<=16'd23725; ROM4[9409]<=16'd57232;
ROM1[9410]<=16'd4771; ROM2[9410]<=16'd0; ROM3[9410]<=16'd23730; ROM4[9410]<=16'd57235;
ROM1[9411]<=16'd4758; ROM2[9411]<=16'd0; ROM3[9411]<=16'd23738; ROM4[9411]<=16'd57235;
ROM1[9412]<=16'd4748; ROM2[9412]<=16'd0; ROM3[9412]<=16'd23728; ROM4[9412]<=16'd57224;
ROM1[9413]<=16'd4770; ROM2[9413]<=16'd0; ROM3[9413]<=16'd23722; ROM4[9413]<=16'd57225;
ROM1[9414]<=16'd4813; ROM2[9414]<=16'd0; ROM3[9414]<=16'd23719; ROM4[9414]<=16'd57231;
ROM1[9415]<=16'd4837; ROM2[9415]<=16'd0; ROM3[9415]<=16'd23717; ROM4[9415]<=16'd57236;
ROM1[9416]<=16'd4836; ROM2[9416]<=16'd0; ROM3[9416]<=16'd23733; ROM4[9416]<=16'd57246;
ROM1[9417]<=16'd4816; ROM2[9417]<=16'd0; ROM3[9417]<=16'd23743; ROM4[9417]<=16'd57246;
ROM1[9418]<=16'd4800; ROM2[9418]<=16'd0; ROM3[9418]<=16'd23753; ROM4[9418]<=16'd57245;
ROM1[9419]<=16'd4792; ROM2[9419]<=16'd0; ROM3[9419]<=16'd23763; ROM4[9419]<=16'd57249;
ROM1[9420]<=16'd4775; ROM2[9420]<=16'd0; ROM3[9420]<=16'd23754; ROM4[9420]<=16'd57243;
ROM1[9421]<=16'd4779; ROM2[9421]<=16'd0; ROM3[9421]<=16'd23740; ROM4[9421]<=16'd57236;
ROM1[9422]<=16'd4804; ROM2[9422]<=16'd0; ROM3[9422]<=16'd23724; ROM4[9422]<=16'd57227;
ROM1[9423]<=16'd4808; ROM2[9423]<=16'd0; ROM3[9423]<=16'd23703; ROM4[9423]<=16'd57213;
ROM1[9424]<=16'd4788; ROM2[9424]<=16'd0; ROM3[9424]<=16'd23694; ROM4[9424]<=16'd57199;
ROM1[9425]<=16'd4775; ROM2[9425]<=16'd0; ROM3[9425]<=16'd23695; ROM4[9425]<=16'd57195;
ROM1[9426]<=16'd4775; ROM2[9426]<=16'd0; ROM3[9426]<=16'd23706; ROM4[9426]<=16'd57204;
ROM1[9427]<=16'd4762; ROM2[9427]<=16'd0; ROM3[9427]<=16'd23709; ROM4[9427]<=16'd57200;
ROM1[9428]<=16'd4741; ROM2[9428]<=16'd0; ROM3[9428]<=16'd23700; ROM4[9428]<=16'd57189;
ROM1[9429]<=16'd4748; ROM2[9429]<=16'd0; ROM3[9429]<=16'd23709; ROM4[9429]<=16'd57197;
ROM1[9430]<=16'd4773; ROM2[9430]<=16'd0; ROM3[9430]<=16'd23710; ROM4[9430]<=16'd57200;
ROM1[9431]<=16'd4792; ROM2[9431]<=16'd0; ROM3[9431]<=16'd23684; ROM4[9431]<=16'd57189;
ROM1[9432]<=16'd4807; ROM2[9432]<=16'd0; ROM3[9432]<=16'd23690; ROM4[9432]<=16'd57200;
ROM1[9433]<=16'd4813; ROM2[9433]<=16'd0; ROM3[9433]<=16'd23710; ROM4[9433]<=16'd57219;
ROM1[9434]<=16'd4805; ROM2[9434]<=16'd0; ROM3[9434]<=16'd23727; ROM4[9434]<=16'd57232;
ROM1[9435]<=16'd4811; ROM2[9435]<=16'd0; ROM3[9435]<=16'd23759; ROM4[9435]<=16'd57257;
ROM1[9436]<=16'd4779; ROM2[9436]<=16'd0; ROM3[9436]<=16'd23744; ROM4[9436]<=16'd57233;
ROM1[9437]<=16'd4741; ROM2[9437]<=16'd0; ROM3[9437]<=16'd23716; ROM4[9437]<=16'd57199;
ROM1[9438]<=16'd4748; ROM2[9438]<=16'd0; ROM3[9438]<=16'd23700; ROM4[9438]<=16'd57191;
ROM1[9439]<=16'd4776; ROM2[9439]<=16'd0; ROM3[9439]<=16'd23680; ROM4[9439]<=16'd57187;
ROM1[9440]<=16'd4794; ROM2[9440]<=16'd0; ROM3[9440]<=16'd23681; ROM4[9440]<=16'd57192;
ROM1[9441]<=16'd4788; ROM2[9441]<=16'd0; ROM3[9441]<=16'd23693; ROM4[9441]<=16'd57200;
ROM1[9442]<=16'd4771; ROM2[9442]<=16'd0; ROM3[9442]<=16'd23707; ROM4[9442]<=16'd57209;
ROM1[9443]<=16'd4763; ROM2[9443]<=16'd0; ROM3[9443]<=16'd23721; ROM4[9443]<=16'd57215;
ROM1[9444]<=16'd4770; ROM2[9444]<=16'd0; ROM3[9444]<=16'd23750; ROM4[9444]<=16'd57239;
ROM1[9445]<=16'd4762; ROM2[9445]<=16'd0; ROM3[9445]<=16'd23747; ROM4[9445]<=16'd57235;
ROM1[9446]<=16'd4748; ROM2[9446]<=16'd0; ROM3[9446]<=16'd23716; ROM4[9446]<=16'd57205;
ROM1[9447]<=16'd4767; ROM2[9447]<=16'd0; ROM3[9447]<=16'd23702; ROM4[9447]<=16'd57198;
ROM1[9448]<=16'd4780; ROM2[9448]<=16'd0; ROM3[9448]<=16'd23683; ROM4[9448]<=16'd57189;
ROM1[9449]<=16'd4788; ROM2[9449]<=16'd0; ROM3[9449]<=16'd23697; ROM4[9449]<=16'd57201;
ROM1[9450]<=16'd4793; ROM2[9450]<=16'd0; ROM3[9450]<=16'd23722; ROM4[9450]<=16'd57219;
ROM1[9451]<=16'd4757; ROM2[9451]<=16'd0; ROM3[9451]<=16'd23707; ROM4[9451]<=16'd57200;
ROM1[9452]<=16'd4716; ROM2[9452]<=16'd0; ROM3[9452]<=16'd23691; ROM4[9452]<=16'd57182;
ROM1[9453]<=16'd4703; ROM2[9453]<=16'd0; ROM3[9453]<=16'd23692; ROM4[9453]<=16'd57181;
ROM1[9454]<=16'd4720; ROM2[9454]<=16'd0; ROM3[9454]<=16'd23696; ROM4[9454]<=16'd57188;
ROM1[9455]<=16'd4756; ROM2[9455]<=16'd0; ROM3[9455]<=16'd23692; ROM4[9455]<=16'd57198;
ROM1[9456]<=16'd4799; ROM2[9456]<=16'd0; ROM3[9456]<=16'd23690; ROM4[9456]<=16'd57205;
ROM1[9457]<=16'd4801; ROM2[9457]<=16'd0; ROM3[9457]<=16'd23684; ROM4[9457]<=16'd57203;
ROM1[9458]<=16'd4786; ROM2[9458]<=16'd0; ROM3[9458]<=16'd23692; ROM4[9458]<=16'd57208;
ROM1[9459]<=16'd4780; ROM2[9459]<=16'd0; ROM3[9459]<=16'd23708; ROM4[9459]<=16'd57217;
ROM1[9460]<=16'd4758; ROM2[9460]<=16'd0; ROM3[9460]<=16'd23700; ROM4[9460]<=16'd57205;
ROM1[9461]<=16'd4732; ROM2[9461]<=16'd0; ROM3[9461]<=16'd23693; ROM4[9461]<=16'd57194;
ROM1[9462]<=16'd4728; ROM2[9462]<=16'd0; ROM3[9462]<=16'd23692; ROM4[9462]<=16'd57192;
ROM1[9463]<=16'd4743; ROM2[9463]<=16'd0; ROM3[9463]<=16'd23686; ROM4[9463]<=16'd57189;
ROM1[9464]<=16'd4782; ROM2[9464]<=16'd0; ROM3[9464]<=16'd23681; ROM4[9464]<=16'd57199;
ROM1[9465]<=16'd4821; ROM2[9465]<=16'd0; ROM3[9465]<=16'd23699; ROM4[9465]<=16'd57222;
ROM1[9466]<=16'd4811; ROM2[9466]<=16'd0; ROM3[9466]<=16'd23708; ROM4[9466]<=16'd57222;
ROM1[9467]<=16'd4774; ROM2[9467]<=16'd0; ROM3[9467]<=16'd23697; ROM4[9467]<=16'd57202;
ROM1[9468]<=16'd4763; ROM2[9468]<=16'd0; ROM3[9468]<=16'd23705; ROM4[9468]<=16'd57206;
ROM1[9469]<=16'd4741; ROM2[9469]<=16'd0; ROM3[9469]<=16'd23705; ROM4[9469]<=16'd57203;
ROM1[9470]<=16'd4727; ROM2[9470]<=16'd0; ROM3[9470]<=16'd23698; ROM4[9470]<=16'd57194;
ROM1[9471]<=16'd4742; ROM2[9471]<=16'd0; ROM3[9471]<=16'd23697; ROM4[9471]<=16'd57198;
ROM1[9472]<=16'd4773; ROM2[9472]<=16'd0; ROM3[9472]<=16'd23695; ROM4[9472]<=16'd57201;
ROM1[9473]<=16'd4804; ROM2[9473]<=16'd0; ROM3[9473]<=16'd23699; ROM4[9473]<=16'd57214;
ROM1[9474]<=16'd4817; ROM2[9474]<=16'd0; ROM3[9474]<=16'd23718; ROM4[9474]<=16'd57234;
ROM1[9475]<=16'd4797; ROM2[9475]<=16'd0; ROM3[9475]<=16'd23721; ROM4[9475]<=16'd57231;
ROM1[9476]<=16'd4786; ROM2[9476]<=16'd0; ROM3[9476]<=16'd23733; ROM4[9476]<=16'd57233;
ROM1[9477]<=16'd4777; ROM2[9477]<=16'd0; ROM3[9477]<=16'd23742; ROM4[9477]<=16'd57230;
ROM1[9478]<=16'd4747; ROM2[9478]<=16'd0; ROM3[9478]<=16'd23725; ROM4[9478]<=16'd57213;
ROM1[9479]<=16'd4766; ROM2[9479]<=16'd0; ROM3[9479]<=16'd23741; ROM4[9479]<=16'd57230;
ROM1[9480]<=16'd4788; ROM2[9480]<=16'd0; ROM3[9480]<=16'd23733; ROM4[9480]<=16'd57225;
ROM1[9481]<=16'd4796; ROM2[9481]<=16'd0; ROM3[9481]<=16'd23700; ROM4[9481]<=16'd57203;
ROM1[9482]<=16'd4798; ROM2[9482]<=16'd0; ROM3[9482]<=16'd23699; ROM4[9482]<=16'd57199;
ROM1[9483]<=16'd4783; ROM2[9483]<=16'd0; ROM3[9483]<=16'd23707; ROM4[9483]<=16'd57198;
ROM1[9484]<=16'd4775; ROM2[9484]<=16'd0; ROM3[9484]<=16'd23723; ROM4[9484]<=16'd57206;
ROM1[9485]<=16'd4770; ROM2[9485]<=16'd0; ROM3[9485]<=16'd23736; ROM4[9485]<=16'd57214;
ROM1[9486]<=16'd4755; ROM2[9486]<=16'd0; ROM3[9486]<=16'd23741; ROM4[9486]<=16'd57218;
ROM1[9487]<=16'd4753; ROM2[9487]<=16'd0; ROM3[9487]<=16'd23742; ROM4[9487]<=16'd57219;
ROM1[9488]<=16'd4768; ROM2[9488]<=16'd0; ROM3[9488]<=16'd23735; ROM4[9488]<=16'd57218;
ROM1[9489]<=16'd4798; ROM2[9489]<=16'd0; ROM3[9489]<=16'd23727; ROM4[9489]<=16'd57220;
ROM1[9490]<=16'd4813; ROM2[9490]<=16'd0; ROM3[9490]<=16'd23725; ROM4[9490]<=16'd57225;
ROM1[9491]<=16'd4799; ROM2[9491]<=16'd0; ROM3[9491]<=16'd23730; ROM4[9491]<=16'd57227;
ROM1[9492]<=16'd4780; ROM2[9492]<=16'd0; ROM3[9492]<=16'd23736; ROM4[9492]<=16'd57229;
ROM1[9493]<=16'd4770; ROM2[9493]<=16'd0; ROM3[9493]<=16'd23749; ROM4[9493]<=16'd57237;
ROM1[9494]<=16'd4760; ROM2[9494]<=16'd0; ROM3[9494]<=16'd23759; ROM4[9494]<=16'd57241;
ROM1[9495]<=16'd4754; ROM2[9495]<=16'd0; ROM3[9495]<=16'd23758; ROM4[9495]<=16'd57235;
ROM1[9496]<=16'd4773; ROM2[9496]<=16'd0; ROM3[9496]<=16'd23758; ROM4[9496]<=16'd57239;
ROM1[9497]<=16'd4812; ROM2[9497]<=16'd0; ROM3[9497]<=16'd23750; ROM4[9497]<=16'd57243;
ROM1[9498]<=16'd4827; ROM2[9498]<=16'd0; ROM3[9498]<=16'd23731; ROM4[9498]<=16'd57230;
ROM1[9499]<=16'd4809; ROM2[9499]<=16'd0; ROM3[9499]<=16'd23720; ROM4[9499]<=16'd57217;
ROM1[9500]<=16'd4780; ROM2[9500]<=16'd0; ROM3[9500]<=16'd23716; ROM4[9500]<=16'd57211;
ROM1[9501]<=16'd4755; ROM2[9501]<=16'd0; ROM3[9501]<=16'd23713; ROM4[9501]<=16'd57201;
ROM1[9502]<=16'd4755; ROM2[9502]<=16'd0; ROM3[9502]<=16'd23725; ROM4[9502]<=16'd57211;
ROM1[9503]<=16'd4755; ROM2[9503]<=16'd0; ROM3[9503]<=16'd23734; ROM4[9503]<=16'd57219;
ROM1[9504]<=16'd4754; ROM2[9504]<=16'd0; ROM3[9504]<=16'd23718; ROM4[9504]<=16'd57209;
ROM1[9505]<=16'd4772; ROM2[9505]<=16'd0; ROM3[9505]<=16'd23702; ROM4[9505]<=16'd57201;
ROM1[9506]<=16'd4796; ROM2[9506]<=16'd0; ROM3[9506]<=16'd23684; ROM4[9506]<=16'd57192;
ROM1[9507]<=16'd4808; ROM2[9507]<=16'd0; ROM3[9507]<=16'd23693; ROM4[9507]<=16'd57204;
ROM1[9508]<=16'd4812; ROM2[9508]<=16'd0; ROM3[9508]<=16'd23718; ROM4[9508]<=16'd57222;
ROM1[9509]<=16'd4799; ROM2[9509]<=16'd0; ROM3[9509]<=16'd23728; ROM4[9509]<=16'd57228;
ROM1[9510]<=16'd4789; ROM2[9510]<=16'd0; ROM3[9510]<=16'd23736; ROM4[9510]<=16'd57238;
ROM1[9511]<=16'd4761; ROM2[9511]<=16'd0; ROM3[9511]<=16'd23728; ROM4[9511]<=16'd57225;
ROM1[9512]<=16'd4732; ROM2[9512]<=16'd0; ROM3[9512]<=16'd23702; ROM4[9512]<=16'd57195;
ROM1[9513]<=16'd4751; ROM2[9513]<=16'd0; ROM3[9513]<=16'd23696; ROM4[9513]<=16'd57195;
ROM1[9514]<=16'd4785; ROM2[9514]<=16'd0; ROM3[9514]<=16'd23688; ROM4[9514]<=16'd57197;
ROM1[9515]<=16'd4802; ROM2[9515]<=16'd0; ROM3[9515]<=16'd23687; ROM4[9515]<=16'd57204;
ROM1[9516]<=16'd4792; ROM2[9516]<=16'd0; ROM3[9516]<=16'd23694; ROM4[9516]<=16'd57205;
ROM1[9517]<=16'd4763; ROM2[9517]<=16'd0; ROM3[9517]<=16'd23692; ROM4[9517]<=16'd57192;
ROM1[9518]<=16'd4737; ROM2[9518]<=16'd0; ROM3[9518]<=16'd23691; ROM4[9518]<=16'd57182;
ROM1[9519]<=16'd4717; ROM2[9519]<=16'd0; ROM3[9519]<=16'd23691; ROM4[9519]<=16'd57175;
ROM1[9520]<=16'd4715; ROM2[9520]<=16'd0; ROM3[9520]<=16'd23698; ROM4[9520]<=16'd57182;
ROM1[9521]<=16'd4735; ROM2[9521]<=16'd0; ROM3[9521]<=16'd23703; ROM4[9521]<=16'd57188;
ROM1[9522]<=16'd4764; ROM2[9522]<=16'd0; ROM3[9522]<=16'd23695; ROM4[9522]<=16'd57185;
ROM1[9523]<=16'd4780; ROM2[9523]<=16'd0; ROM3[9523]<=16'd23683; ROM4[9523]<=16'd57179;
ROM1[9524]<=16'd4778; ROM2[9524]<=16'd0; ROM3[9524]<=16'd23689; ROM4[9524]<=16'd57184;
ROM1[9525]<=16'd4765; ROM2[9525]<=16'd0; ROM3[9525]<=16'd23701; ROM4[9525]<=16'd57192;
ROM1[9526]<=16'd4752; ROM2[9526]<=16'd0; ROM3[9526]<=16'd23712; ROM4[9526]<=16'd57194;
ROM1[9527]<=16'd4744; ROM2[9527]<=16'd0; ROM3[9527]<=16'd23723; ROM4[9527]<=16'd57203;
ROM1[9528]<=16'd4738; ROM2[9528]<=16'd0; ROM3[9528]<=16'd23732; ROM4[9528]<=16'd57208;
ROM1[9529]<=16'd4748; ROM2[9529]<=16'd0; ROM3[9529]<=16'd23728; ROM4[9529]<=16'd57204;
ROM1[9530]<=16'd4772; ROM2[9530]<=16'd0; ROM3[9530]<=16'd23718; ROM4[9530]<=16'd57204;
ROM1[9531]<=16'd4808; ROM2[9531]<=16'd0; ROM3[9531]<=16'd23713; ROM4[9531]<=16'd57209;
ROM1[9532]<=16'd4815; ROM2[9532]<=16'd0; ROM3[9532]<=16'd23716; ROM4[9532]<=16'd57210;
ROM1[9533]<=16'd4810; ROM2[9533]<=16'd0; ROM3[9533]<=16'd23739; ROM4[9533]<=16'd57227;
ROM1[9534]<=16'd4805; ROM2[9534]<=16'd0; ROM3[9534]<=16'd23759; ROM4[9534]<=16'd57243;
ROM1[9535]<=16'd4794; ROM2[9535]<=16'd0; ROM3[9535]<=16'd23762; ROM4[9535]<=16'd57243;
ROM1[9536]<=16'd4762; ROM2[9536]<=16'd0; ROM3[9536]<=16'd23750; ROM4[9536]<=16'd57225;
ROM1[9537]<=16'd4739; ROM2[9537]<=16'd0; ROM3[9537]<=16'd23735; ROM4[9537]<=16'd57205;
ROM1[9538]<=16'd4758; ROM2[9538]<=16'd0; ROM3[9538]<=16'd23740; ROM4[9538]<=16'd57209;
ROM1[9539]<=16'd4805; ROM2[9539]<=16'd0; ROM3[9539]<=16'd23754; ROM4[9539]<=16'd57231;
ROM1[9540]<=16'd4824; ROM2[9540]<=16'd0; ROM3[9540]<=16'd23761; ROM4[9540]<=16'd57245;
ROM1[9541]<=16'd4811; ROM2[9541]<=16'd0; ROM3[9541]<=16'd23769; ROM4[9541]<=16'd57250;
ROM1[9542]<=16'd4801; ROM2[9542]<=16'd0; ROM3[9542]<=16'd23786; ROM4[9542]<=16'd57257;
ROM1[9543]<=16'd4784; ROM2[9543]<=16'd0; ROM3[9543]<=16'd23783; ROM4[9543]<=16'd57252;
ROM1[9544]<=16'd4780; ROM2[9544]<=16'd0; ROM3[9544]<=16'd23796; ROM4[9544]<=16'd57267;
ROM1[9545]<=16'd4789; ROM2[9545]<=16'd0; ROM3[9545]<=16'd23813; ROM4[9545]<=16'd57283;
ROM1[9546]<=16'd4777; ROM2[9546]<=16'd0; ROM3[9546]<=16'd23782; ROM4[9546]<=16'd57258;
ROM1[9547]<=16'd4790; ROM2[9547]<=16'd0; ROM3[9547]<=16'd23753; ROM4[9547]<=16'd57235;
ROM1[9548]<=16'd4820; ROM2[9548]<=16'd0; ROM3[9548]<=16'd23745; ROM4[9548]<=16'd57233;
ROM1[9549]<=16'd4815; ROM2[9549]<=16'd0; ROM3[9549]<=16'd23741; ROM4[9549]<=16'd57229;
ROM1[9550]<=16'd4809; ROM2[9550]<=16'd0; ROM3[9550]<=16'd23754; ROM4[9550]<=16'd57240;
ROM1[9551]<=16'd4799; ROM2[9551]<=16'd0; ROM3[9551]<=16'd23763; ROM4[9551]<=16'd57244;
ROM1[9552]<=16'd4782; ROM2[9552]<=16'd0; ROM3[9552]<=16'd23758; ROM4[9552]<=16'd57237;
ROM1[9553]<=16'd4773; ROM2[9553]<=16'd0; ROM3[9553]<=16'd23753; ROM4[9553]<=16'd57233;
ROM1[9554]<=16'd4774; ROM2[9554]<=16'd0; ROM3[9554]<=16'd23748; ROM4[9554]<=16'd57226;
ROM1[9555]<=16'd4805; ROM2[9555]<=16'd0; ROM3[9555]<=16'd23745; ROM4[9555]<=16'd57228;
ROM1[9556]<=16'd4835; ROM2[9556]<=16'd0; ROM3[9556]<=16'd23735; ROM4[9556]<=16'd57226;
ROM1[9557]<=16'd4835; ROM2[9557]<=16'd0; ROM3[9557]<=16'd23733; ROM4[9557]<=16'd57227;
ROM1[9558]<=16'd4826; ROM2[9558]<=16'd0; ROM3[9558]<=16'd23743; ROM4[9558]<=16'd57236;
ROM1[9559]<=16'd4807; ROM2[9559]<=16'd0; ROM3[9559]<=16'd23748; ROM4[9559]<=16'd57235;
ROM1[9560]<=16'd4791; ROM2[9560]<=16'd0; ROM3[9560]<=16'd23750; ROM4[9560]<=16'd57234;
ROM1[9561]<=16'd4770; ROM2[9561]<=16'd0; ROM3[9561]<=16'd23749; ROM4[9561]<=16'd57227;
ROM1[9562]<=16'd4765; ROM2[9562]<=16'd0; ROM3[9562]<=16'd23743; ROM4[9562]<=16'd57221;
ROM1[9563]<=16'd4782; ROM2[9563]<=16'd0; ROM3[9563]<=16'd23733; ROM4[9563]<=16'd57224;
ROM1[9564]<=16'd4814; ROM2[9564]<=16'd0; ROM3[9564]<=16'd23727; ROM4[9564]<=16'd57227;
ROM1[9565]<=16'd4828; ROM2[9565]<=16'd0; ROM3[9565]<=16'd23723; ROM4[9565]<=16'd57230;
ROM1[9566]<=16'd4817; ROM2[9566]<=16'd0; ROM3[9566]<=16'd23728; ROM4[9566]<=16'd57234;
ROM1[9567]<=16'd4805; ROM2[9567]<=16'd0; ROM3[9567]<=16'd23739; ROM4[9567]<=16'd57245;
ROM1[9568]<=16'd4800; ROM2[9568]<=16'd0; ROM3[9568]<=16'd23754; ROM4[9568]<=16'd57257;
ROM1[9569]<=16'd4785; ROM2[9569]<=16'd0; ROM3[9569]<=16'd23760; ROM4[9569]<=16'd57257;
ROM1[9570]<=16'd4783; ROM2[9570]<=16'd0; ROM3[9570]<=16'd23764; ROM4[9570]<=16'd57259;
ROM1[9571]<=16'd4793; ROM2[9571]<=16'd0; ROM3[9571]<=16'd23759; ROM4[9571]<=16'd57254;
ROM1[9572]<=16'd4800; ROM2[9572]<=16'd0; ROM3[9572]<=16'd23727; ROM4[9572]<=16'd57231;
ROM1[9573]<=16'd4815; ROM2[9573]<=16'd0; ROM3[9573]<=16'd23708; ROM4[9573]<=16'd57224;
ROM1[9574]<=16'd4802; ROM2[9574]<=16'd0; ROM3[9574]<=16'd23702; ROM4[9574]<=16'd57214;
ROM1[9575]<=16'd4764; ROM2[9575]<=16'd0; ROM3[9575]<=16'd23689; ROM4[9575]<=16'd57191;
ROM1[9576]<=16'd4742; ROM2[9576]<=16'd0; ROM3[9576]<=16'd23691; ROM4[9576]<=16'd57181;
ROM1[9577]<=16'd4733; ROM2[9577]<=16'd0; ROM3[9577]<=16'd23701; ROM4[9577]<=16'd57180;
ROM1[9578]<=16'd4724; ROM2[9578]<=16'd0; ROM3[9578]<=16'd23704; ROM4[9578]<=16'd57180;
ROM1[9579]<=16'd4740; ROM2[9579]<=16'd0; ROM3[9579]<=16'd23712; ROM4[9579]<=16'd57188;
ROM1[9580]<=16'd4770; ROM2[9580]<=16'd0; ROM3[9580]<=16'd23709; ROM4[9580]<=16'd57190;
ROM1[9581]<=16'd4796; ROM2[9581]<=16'd0; ROM3[9581]<=16'd23695; ROM4[9581]<=16'd57186;
ROM1[9582]<=16'd4805; ROM2[9582]<=16'd0; ROM3[9582]<=16'd23706; ROM4[9582]<=16'd57194;
ROM1[9583]<=16'd4801; ROM2[9583]<=16'd0; ROM3[9583]<=16'd23726; ROM4[9583]<=16'd57207;
ROM1[9584]<=16'd4760; ROM2[9584]<=16'd0; ROM3[9584]<=16'd23712; ROM4[9584]<=16'd57186;
ROM1[9585]<=16'd4728; ROM2[9585]<=16'd0; ROM3[9585]<=16'd23699; ROM4[9585]<=16'd57166;
ROM1[9586]<=16'd4709; ROM2[9586]<=16'd0; ROM3[9586]<=16'd23696; ROM4[9586]<=16'd57161;
ROM1[9587]<=16'd4705; ROM2[9587]<=16'd0; ROM3[9587]<=16'd23693; ROM4[9587]<=16'd57155;
ROM1[9588]<=16'd4742; ROM2[9588]<=16'd0; ROM3[9588]<=16'd23707; ROM4[9588]<=16'd57171;
ROM1[9589]<=16'd4783; ROM2[9589]<=16'd0; ROM3[9589]<=16'd23706; ROM4[9589]<=16'd57186;
ROM1[9590]<=16'd4791; ROM2[9590]<=16'd0; ROM3[9590]<=16'd23699; ROM4[9590]<=16'd57185;
ROM1[9591]<=16'd4775; ROM2[9591]<=16'd0; ROM3[9591]<=16'd23708; ROM4[9591]<=16'd57192;
ROM1[9592]<=16'd4770; ROM2[9592]<=16'd0; ROM3[9592]<=16'd23725; ROM4[9592]<=16'd57208;
ROM1[9593]<=16'd4769; ROM2[9593]<=16'd0; ROM3[9593]<=16'd23747; ROM4[9593]<=16'd57224;
ROM1[9594]<=16'd4760; ROM2[9594]<=16'd0; ROM3[9594]<=16'd23768; ROM4[9594]<=16'd57236;
ROM1[9595]<=16'd4760; ROM2[9595]<=16'd0; ROM3[9595]<=16'd23776; ROM4[9595]<=16'd57242;
ROM1[9596]<=16'd4774; ROM2[9596]<=16'd0; ROM3[9596]<=16'd23777; ROM4[9596]<=16'd57247;
ROM1[9597]<=16'd4805; ROM2[9597]<=16'd0; ROM3[9597]<=16'd23774; ROM4[9597]<=16'd57254;
ROM1[9598]<=16'd4831; ROM2[9598]<=16'd0; ROM3[9598]<=16'd23772; ROM4[9598]<=16'd57260;
ROM1[9599]<=16'd4830; ROM2[9599]<=16'd0; ROM3[9599]<=16'd23780; ROM4[9599]<=16'd57267;
ROM1[9600]<=16'd4819; ROM2[9600]<=16'd0; ROM3[9600]<=16'd23797; ROM4[9600]<=16'd57277;
ROM1[9601]<=16'd4810; ROM2[9601]<=16'd0; ROM3[9601]<=16'd23812; ROM4[9601]<=16'd57281;
ROM1[9602]<=16'd4801; ROM2[9602]<=16'd0; ROM3[9602]<=16'd23819; ROM4[9602]<=16'd57284;
ROM1[9603]<=16'd4785; ROM2[9603]<=16'd0; ROM3[9603]<=16'd23817; ROM4[9603]<=16'd57274;
ROM1[9604]<=16'd4794; ROM2[9604]<=16'd0; ROM3[9604]<=16'd23821; ROM4[9604]<=16'd57276;
ROM1[9605]<=16'd4812; ROM2[9605]<=16'd0; ROM3[9605]<=16'd23796; ROM4[9605]<=16'd57264;
ROM1[9606]<=16'd4822; ROM2[9606]<=16'd0; ROM3[9606]<=16'd23757; ROM4[9606]<=16'd57237;
ROM1[9607]<=16'd4824; ROM2[9607]<=16'd0; ROM3[9607]<=16'd23747; ROM4[9607]<=16'd57234;
ROM1[9608]<=16'd4808; ROM2[9608]<=16'd0; ROM3[9608]<=16'd23747; ROM4[9608]<=16'd57229;
ROM1[9609]<=16'd4804; ROM2[9609]<=16'd0; ROM3[9609]<=16'd23762; ROM4[9609]<=16'd57237;
ROM1[9610]<=16'd4815; ROM2[9610]<=16'd0; ROM3[9610]<=16'd23783; ROM4[9610]<=16'd57250;
ROM1[9611]<=16'd4793; ROM2[9611]<=16'd0; ROM3[9611]<=16'd23777; ROM4[9611]<=16'd57234;
ROM1[9612]<=16'd4771; ROM2[9612]<=16'd0; ROM3[9612]<=16'd23750; ROM4[9612]<=16'd57211;
ROM1[9613]<=16'd4783; ROM2[9613]<=16'd0; ROM3[9613]<=16'd23728; ROM4[9613]<=16'd57198;
ROM1[9614]<=16'd4807; ROM2[9614]<=16'd0; ROM3[9614]<=16'd23707; ROM4[9614]<=16'd57187;
ROM1[9615]<=16'd4822; ROM2[9615]<=16'd0; ROM3[9615]<=16'd23698; ROM4[9615]<=16'd57187;
ROM1[9616]<=16'd4819; ROM2[9616]<=16'd0; ROM3[9616]<=16'd23706; ROM4[9616]<=16'd57193;
ROM1[9617]<=16'd4809; ROM2[9617]<=16'd0; ROM3[9617]<=16'd23729; ROM4[9617]<=16'd57202;
ROM1[9618]<=16'd4785; ROM2[9618]<=16'd0; ROM3[9618]<=16'd23724; ROM4[9618]<=16'd57192;
ROM1[9619]<=16'd4760; ROM2[9619]<=16'd0; ROM3[9619]<=16'd23719; ROM4[9619]<=16'd57184;
ROM1[9620]<=16'd4759; ROM2[9620]<=16'd0; ROM3[9620]<=16'd23727; ROM4[9620]<=16'd57191;
ROM1[9621]<=16'd4761; ROM2[9621]<=16'd0; ROM3[9621]<=16'd23704; ROM4[9621]<=16'd57174;
ROM1[9622]<=16'd4782; ROM2[9622]<=16'd0; ROM3[9622]<=16'd23684; ROM4[9622]<=16'd57169;
ROM1[9623]<=16'd4807; ROM2[9623]<=16'd0; ROM3[9623]<=16'd23678; ROM4[9623]<=16'd57178;
ROM1[9624]<=16'd4803; ROM2[9624]<=16'd0; ROM3[9624]<=16'd23680; ROM4[9624]<=16'd57178;
ROM1[9625]<=16'd4776; ROM2[9625]<=16'd0; ROM3[9625]<=16'd23682; ROM4[9625]<=16'd57175;
ROM1[9626]<=16'd4762; ROM2[9626]<=16'd0; ROM3[9626]<=16'd23697; ROM4[9626]<=16'd57186;
ROM1[9627]<=16'd4757; ROM2[9627]<=16'd0; ROM3[9627]<=16'd23716; ROM4[9627]<=16'd57196;
ROM1[9628]<=16'd4745; ROM2[9628]<=16'd0; ROM3[9628]<=16'd23717; ROM4[9628]<=16'd57195;
ROM1[9629]<=16'd4752; ROM2[9629]<=16'd0; ROM3[9629]<=16'd23719; ROM4[9629]<=16'd57200;
ROM1[9630]<=16'd4783; ROM2[9630]<=16'd0; ROM3[9630]<=16'd23720; ROM4[9630]<=16'd57202;
ROM1[9631]<=16'd4818; ROM2[9631]<=16'd0; ROM3[9631]<=16'd23716; ROM4[9631]<=16'd57208;
ROM1[9632]<=16'd4822; ROM2[9632]<=16'd0; ROM3[9632]<=16'd23720; ROM4[9632]<=16'd57214;
ROM1[9633]<=16'd4812; ROM2[9633]<=16'd0; ROM3[9633]<=16'd23739; ROM4[9633]<=16'd57223;
ROM1[9634]<=16'd4800; ROM2[9634]<=16'd0; ROM3[9634]<=16'd23757; ROM4[9634]<=16'd57232;
ROM1[9635]<=16'd4789; ROM2[9635]<=16'd0; ROM3[9635]<=16'd23763; ROM4[9635]<=16'd57233;
ROM1[9636]<=16'd4777; ROM2[9636]<=16'd0; ROM3[9636]<=16'd23776; ROM4[9636]<=16'd57235;
ROM1[9637]<=16'd4782; ROM2[9637]<=16'd0; ROM3[9637]<=16'd23780; ROM4[9637]<=16'd57240;
ROM1[9638]<=16'd4809; ROM2[9638]<=16'd0; ROM3[9638]<=16'd23780; ROM4[9638]<=16'd57246;
ROM1[9639]<=16'd4844; ROM2[9639]<=16'd0; ROM3[9639]<=16'd23772; ROM4[9639]<=16'd57246;
ROM1[9640]<=16'd4860; ROM2[9640]<=16'd0; ROM3[9640]<=16'd23772; ROM4[9640]<=16'd57247;
ROM1[9641]<=16'd4862; ROM2[9641]<=16'd0; ROM3[9641]<=16'd23790; ROM4[9641]<=16'd57261;
ROM1[9642]<=16'd4828; ROM2[9642]<=16'd0; ROM3[9642]<=16'd23782; ROM4[9642]<=16'd57247;
ROM1[9643]<=16'd4800; ROM2[9643]<=16'd0; ROM3[9643]<=16'd23772; ROM4[9643]<=16'd57228;
ROM1[9644]<=16'd4804; ROM2[9644]<=16'd0; ROM3[9644]<=16'd23794; ROM4[9644]<=16'd57244;
ROM1[9645]<=16'd4791; ROM2[9645]<=16'd0; ROM3[9645]<=16'd23791; ROM4[9645]<=16'd57237;
ROM1[9646]<=16'd4797; ROM2[9646]<=16'd0; ROM3[9646]<=16'd23779; ROM4[9646]<=16'd57230;
ROM1[9647]<=16'd4819; ROM2[9647]<=16'd0; ROM3[9647]<=16'd23764; ROM4[9647]<=16'd57227;
ROM1[9648]<=16'd4815; ROM2[9648]<=16'd0; ROM3[9648]<=16'd23729; ROM4[9648]<=16'd57200;
ROM1[9649]<=16'd4799; ROM2[9649]<=16'd0; ROM3[9649]<=16'd23718; ROM4[9649]<=16'd57193;
ROM1[9650]<=16'd4789; ROM2[9650]<=16'd0; ROM3[9650]<=16'd23734; ROM4[9650]<=16'd57203;
ROM1[9651]<=16'd4784; ROM2[9651]<=16'd0; ROM3[9651]<=16'd23749; ROM4[9651]<=16'd57214;
ROM1[9652]<=16'd4779; ROM2[9652]<=16'd0; ROM3[9652]<=16'd23757; ROM4[9652]<=16'd57220;
ROM1[9653]<=16'd4771; ROM2[9653]<=16'd0; ROM3[9653]<=16'd23762; ROM4[9653]<=16'd57218;
ROM1[9654]<=16'd4792; ROM2[9654]<=16'd0; ROM3[9654]<=16'd23773; ROM4[9654]<=16'd57230;
ROM1[9655]<=16'd4833; ROM2[9655]<=16'd0; ROM3[9655]<=16'd23779; ROM4[9655]<=16'd57244;
ROM1[9656]<=16'd4845; ROM2[9656]<=16'd0; ROM3[9656]<=16'd23747; ROM4[9656]<=16'd57228;
ROM1[9657]<=16'd4830; ROM2[9657]<=16'd0; ROM3[9657]<=16'd23718; ROM4[9657]<=16'd57205;
ROM1[9658]<=16'd4805; ROM2[9658]<=16'd0; ROM3[9658]<=16'd23704; ROM4[9658]<=16'd57190;
ROM1[9659]<=16'd4782; ROM2[9659]<=16'd0; ROM3[9659]<=16'd23703; ROM4[9659]<=16'd57184;
ROM1[9660]<=16'd4772; ROM2[9660]<=16'd0; ROM3[9660]<=16'd23713; ROM4[9660]<=16'd57189;
ROM1[9661]<=16'd4759; ROM2[9661]<=16'd0; ROM3[9661]<=16'd23717; ROM4[9661]<=16'd57191;
ROM1[9662]<=16'd4757; ROM2[9662]<=16'd0; ROM3[9662]<=16'd23709; ROM4[9662]<=16'd57185;
ROM1[9663]<=16'd4778; ROM2[9663]<=16'd0; ROM3[9663]<=16'd23697; ROM4[9663]<=16'd57182;
ROM1[9664]<=16'd4814; ROM2[9664]<=16'd0; ROM3[9664]<=16'd23686; ROM4[9664]<=16'd57184;
ROM1[9665]<=16'd4836; ROM2[9665]<=16'd0; ROM3[9665]<=16'd23688; ROM4[9665]<=16'd57194;
ROM1[9666]<=16'd4829; ROM2[9666]<=16'd0; ROM3[9666]<=16'd23696; ROM4[9666]<=16'd57202;
ROM1[9667]<=16'd4815; ROM2[9667]<=16'd0; ROM3[9667]<=16'd23713; ROM4[9667]<=16'd57210;
ROM1[9668]<=16'd4821; ROM2[9668]<=16'd0; ROM3[9668]<=16'd23739; ROM4[9668]<=16'd57229;
ROM1[9669]<=16'd4802; ROM2[9669]<=16'd0; ROM3[9669]<=16'd23742; ROM4[9669]<=16'd57224;
ROM1[9670]<=16'd4776; ROM2[9670]<=16'd0; ROM3[9670]<=16'd23725; ROM4[9670]<=16'd57205;
ROM1[9671]<=16'd4774; ROM2[9671]<=16'd0; ROM3[9671]<=16'd23708; ROM4[9671]<=16'd57189;
ROM1[9672]<=16'd4795; ROM2[9672]<=16'd0; ROM3[9672]<=16'd23693; ROM4[9672]<=16'd57182;
ROM1[9673]<=16'd4828; ROM2[9673]<=16'd0; ROM3[9673]<=16'd23692; ROM4[9673]<=16'd57192;
ROM1[9674]<=16'd4829; ROM2[9674]<=16'd0; ROM3[9674]<=16'd23703; ROM4[9674]<=16'd57199;
ROM1[9675]<=16'd4818; ROM2[9675]<=16'd0; ROM3[9675]<=16'd23723; ROM4[9675]<=16'd57207;
ROM1[9676]<=16'd4795; ROM2[9676]<=16'd0; ROM3[9676]<=16'd23728; ROM4[9676]<=16'd57202;
ROM1[9677]<=16'd4770; ROM2[9677]<=16'd0; ROM3[9677]<=16'd23729; ROM4[9677]<=16'd57192;
ROM1[9678]<=16'd4765; ROM2[9678]<=16'd0; ROM3[9678]<=16'd23743; ROM4[9678]<=16'd57199;
ROM1[9679]<=16'd4775; ROM2[9679]<=16'd0; ROM3[9679]<=16'd23745; ROM4[9679]<=16'd57204;
ROM1[9680]<=16'd4809; ROM2[9680]<=16'd0; ROM3[9680]<=16'd23746; ROM4[9680]<=16'd57214;
ROM1[9681]<=16'd4846; ROM2[9681]<=16'd0; ROM3[9681]<=16'd23742; ROM4[9681]<=16'd57223;
ROM1[9682]<=16'd4851; ROM2[9682]<=16'd0; ROM3[9682]<=16'd23746; ROM4[9682]<=16'd57228;
ROM1[9683]<=16'd4847; ROM2[9683]<=16'd0; ROM3[9683]<=16'd23768; ROM4[9683]<=16'd57246;
ROM1[9684]<=16'd4846; ROM2[9684]<=16'd0; ROM3[9684]<=16'd23791; ROM4[9684]<=16'd57265;
ROM1[9685]<=16'd4816; ROM2[9685]<=16'd0; ROM3[9685]<=16'd23786; ROM4[9685]<=16'd57253;
ROM1[9686]<=16'd4777; ROM2[9686]<=16'd0; ROM3[9686]<=16'd23766; ROM4[9686]<=16'd57230;
ROM1[9687]<=16'd4773; ROM2[9687]<=16'd0; ROM3[9687]<=16'd23759; ROM4[9687]<=16'd57224;
ROM1[9688]<=16'd4787; ROM2[9688]<=16'd0; ROM3[9688]<=16'd23749; ROM4[9688]<=16'd57219;
ROM1[9689]<=16'd4830; ROM2[9689]<=16'd0; ROM3[9689]<=16'd23748; ROM4[9689]<=16'd57229;
ROM1[9690]<=16'd4862; ROM2[9690]<=16'd0; ROM3[9690]<=16'd23761; ROM4[9690]<=16'd57244;
ROM1[9691]<=16'd4859; ROM2[9691]<=16'd0; ROM3[9691]<=16'd23769; ROM4[9691]<=16'd57251;
ROM1[9692]<=16'd4844; ROM2[9692]<=16'd0; ROM3[9692]<=16'd23781; ROM4[9692]<=16'd57259;
ROM1[9693]<=16'd4809; ROM2[9693]<=16'd0; ROM3[9693]<=16'd23772; ROM4[9693]<=16'd57235;
ROM1[9694]<=16'd4763; ROM2[9694]<=16'd0; ROM3[9694]<=16'd23741; ROM4[9694]<=16'd57200;
ROM1[9695]<=16'd4735; ROM2[9695]<=16'd0; ROM3[9695]<=16'd23722; ROM4[9695]<=16'd57178;
ROM1[9696]<=16'd4738; ROM2[9696]<=16'd0; ROM3[9696]<=16'd23709; ROM4[9696]<=16'd57167;
ROM1[9697]<=16'd4788; ROM2[9697]<=16'd0; ROM3[9697]<=16'd23713; ROM4[9697]<=16'd57188;
ROM1[9698]<=16'd4834; ROM2[9698]<=16'd0; ROM3[9698]<=16'd23731; ROM4[9698]<=16'd57211;
ROM1[9699]<=16'd4828; ROM2[9699]<=16'd0; ROM3[9699]<=16'd23733; ROM4[9699]<=16'd57211;
ROM1[9700]<=16'd4804; ROM2[9700]<=16'd0; ROM3[9700]<=16'd23722; ROM4[9700]<=16'd57199;
ROM1[9701]<=16'd4810; ROM2[9701]<=16'd0; ROM3[9701]<=16'd23744; ROM4[9701]<=16'd57220;
ROM1[9702]<=16'd4809; ROM2[9702]<=16'd0; ROM3[9702]<=16'd23769; ROM4[9702]<=16'd57237;
ROM1[9703]<=16'd4781; ROM2[9703]<=16'd0; ROM3[9703]<=16'd23760; ROM4[9703]<=16'd57223;
ROM1[9704]<=16'd4780; ROM2[9704]<=16'd0; ROM3[9704]<=16'd23746; ROM4[9704]<=16'd57213;
ROM1[9705]<=16'd4797; ROM2[9705]<=16'd0; ROM3[9705]<=16'd23727; ROM4[9705]<=16'd57200;
ROM1[9706]<=16'd4823; ROM2[9706]<=16'd0; ROM3[9706]<=16'd23712; ROM4[9706]<=16'd57196;
ROM1[9707]<=16'd4828; ROM2[9707]<=16'd0; ROM3[9707]<=16'd23714; ROM4[9707]<=16'd57202;
ROM1[9708]<=16'd4816; ROM2[9708]<=16'd0; ROM3[9708]<=16'd23727; ROM4[9708]<=16'd57207;
ROM1[9709]<=16'd4801; ROM2[9709]<=16'd0; ROM3[9709]<=16'd23738; ROM4[9709]<=16'd57210;
ROM1[9710]<=16'd4795; ROM2[9710]<=16'd0; ROM3[9710]<=16'd23750; ROM4[9710]<=16'd57221;
ROM1[9711]<=16'd4788; ROM2[9711]<=16'd0; ROM3[9711]<=16'd23758; ROM4[9711]<=16'd57224;
ROM1[9712]<=16'd4795; ROM2[9712]<=16'd0; ROM3[9712]<=16'd23771; ROM4[9712]<=16'd57234;
ROM1[9713]<=16'd4821; ROM2[9713]<=16'd0; ROM3[9713]<=16'd23779; ROM4[9713]<=16'd57248;
ROM1[9714]<=16'd4840; ROM2[9714]<=16'd0; ROM3[9714]<=16'd23750; ROM4[9714]<=16'd57235;
ROM1[9715]<=16'd4841; ROM2[9715]<=16'd0; ROM3[9715]<=16'd23733; ROM4[9715]<=16'd57227;
ROM1[9716]<=16'd4825; ROM2[9716]<=16'd0; ROM3[9716]<=16'd23734; ROM4[9716]<=16'd57221;
ROM1[9717]<=16'd4797; ROM2[9717]<=16'd0; ROM3[9717]<=16'd23733; ROM4[9717]<=16'd57209;
ROM1[9718]<=16'd4786; ROM2[9718]<=16'd0; ROM3[9718]<=16'd23741; ROM4[9718]<=16'd57216;
ROM1[9719]<=16'd4780; ROM2[9719]<=16'd0; ROM3[9719]<=16'd23754; ROM4[9719]<=16'd57226;
ROM1[9720]<=16'd4780; ROM2[9720]<=16'd0; ROM3[9720]<=16'd23752; ROM4[9720]<=16'd57230;
ROM1[9721]<=16'd4798; ROM2[9721]<=16'd0; ROM3[9721]<=16'd23746; ROM4[9721]<=16'd57229;
ROM1[9722]<=16'd4836; ROM2[9722]<=16'd0; ROM3[9722]<=16'd23744; ROM4[9722]<=16'd57233;
ROM1[9723]<=16'd4843; ROM2[9723]<=16'd0; ROM3[9723]<=16'd23720; ROM4[9723]<=16'd57217;
ROM1[9724]<=16'd4814; ROM2[9724]<=16'd0; ROM3[9724]<=16'd23704; ROM4[9724]<=16'd57199;
ROM1[9725]<=16'd4792; ROM2[9725]<=16'd0; ROM3[9725]<=16'd23707; ROM4[9725]<=16'd57199;
ROM1[9726]<=16'd4780; ROM2[9726]<=16'd0; ROM3[9726]<=16'd23718; ROM4[9726]<=16'd57200;
ROM1[9727]<=16'd4798; ROM2[9727]<=16'd0; ROM3[9727]<=16'd23754; ROM4[9727]<=16'd57230;
ROM1[9728]<=16'd4812; ROM2[9728]<=16'd0; ROM3[9728]<=16'd23776; ROM4[9728]<=16'd57255;
ROM1[9729]<=16'd4807; ROM2[9729]<=16'd0; ROM3[9729]<=16'd23756; ROM4[9729]<=16'd57236;
ROM1[9730]<=16'd4825; ROM2[9730]<=16'd0; ROM3[9730]<=16'd23740; ROM4[9730]<=16'd57228;
ROM1[9731]<=16'd4862; ROM2[9731]<=16'd0; ROM3[9731]<=16'd23738; ROM4[9731]<=16'd57240;
ROM1[9732]<=16'd4854; ROM2[9732]<=16'd0; ROM3[9732]<=16'd23733; ROM4[9732]<=16'd57232;
ROM1[9733]<=16'd4829; ROM2[9733]<=16'd0; ROM3[9733]<=16'd23730; ROM4[9733]<=16'd57224;
ROM1[9734]<=16'd4807; ROM2[9734]<=16'd0; ROM3[9734]<=16'd23732; ROM4[9734]<=16'd57223;
ROM1[9735]<=16'd4791; ROM2[9735]<=16'd0; ROM3[9735]<=16'd23734; ROM4[9735]<=16'd57216;
ROM1[9736]<=16'd4779; ROM2[9736]<=16'd0; ROM3[9736]<=16'd23730; ROM4[9736]<=16'd57215;
ROM1[9737]<=16'd4788; ROM2[9737]<=16'd0; ROM3[9737]<=16'd23737; ROM4[9737]<=16'd57222;
ROM1[9738]<=16'd4812; ROM2[9738]<=16'd0; ROM3[9738]<=16'd23735; ROM4[9738]<=16'd57225;
ROM1[9739]<=16'd4839; ROM2[9739]<=16'd0; ROM3[9739]<=16'd23720; ROM4[9739]<=16'd57221;
ROM1[9740]<=16'd4853; ROM2[9740]<=16'd0; ROM3[9740]<=16'd23718; ROM4[9740]<=16'd57221;
ROM1[9741]<=16'd4839; ROM2[9741]<=16'd0; ROM3[9741]<=16'd23726; ROM4[9741]<=16'd57227;
ROM1[9742]<=16'd4825; ROM2[9742]<=16'd0; ROM3[9742]<=16'd23740; ROM4[9742]<=16'd57229;
ROM1[9743]<=16'd4823; ROM2[9743]<=16'd0; ROM3[9743]<=16'd23755; ROM4[9743]<=16'd57238;
ROM1[9744]<=16'd4800; ROM2[9744]<=16'd0; ROM3[9744]<=16'd23754; ROM4[9744]<=16'd57234;
ROM1[9745]<=16'd4781; ROM2[9745]<=16'd0; ROM3[9745]<=16'd23745; ROM4[9745]<=16'd57225;
ROM1[9746]<=16'd4788; ROM2[9746]<=16'd0; ROM3[9746]<=16'd23734; ROM4[9746]<=16'd57222;
ROM1[9747]<=16'd4810; ROM2[9747]<=16'd0; ROM3[9747]<=16'd23716; ROM4[9747]<=16'd57212;
ROM1[9748]<=16'd4831; ROM2[9748]<=16'd0; ROM3[9748]<=16'd23717; ROM4[9748]<=16'd57216;
ROM1[9749]<=16'd4826; ROM2[9749]<=16'd0; ROM3[9749]<=16'd23727; ROM4[9749]<=16'd57222;
ROM1[9750]<=16'd4808; ROM2[9750]<=16'd0; ROM3[9750]<=16'd23735; ROM4[9750]<=16'd57222;
ROM1[9751]<=16'd4793; ROM2[9751]<=16'd0; ROM3[9751]<=16'd23739; ROM4[9751]<=16'd57219;
ROM1[9752]<=16'd4784; ROM2[9752]<=16'd0; ROM3[9752]<=16'd23744; ROM4[9752]<=16'd57222;
ROM1[9753]<=16'd4781; ROM2[9753]<=16'd0; ROM3[9753]<=16'd23757; ROM4[9753]<=16'd57229;
ROM1[9754]<=16'd4784; ROM2[9754]<=16'd0; ROM3[9754]<=16'd23761; ROM4[9754]<=16'd57230;
ROM1[9755]<=16'd4798; ROM2[9755]<=16'd0; ROM3[9755]<=16'd23746; ROM4[9755]<=16'd57226;
ROM1[9756]<=16'd4823; ROM2[9756]<=16'd0; ROM3[9756]<=16'd23728; ROM4[9756]<=16'd57220;
ROM1[9757]<=16'd4836; ROM2[9757]<=16'd0; ROM3[9757]<=16'd23729; ROM4[9757]<=16'd57223;
ROM1[9758]<=16'd4828; ROM2[9758]<=16'd0; ROM3[9758]<=16'd23736; ROM4[9758]<=16'd57228;
ROM1[9759]<=16'd4804; ROM2[9759]<=16'd0; ROM3[9759]<=16'd23744; ROM4[9759]<=16'd57226;
ROM1[9760]<=16'd4789; ROM2[9760]<=16'd0; ROM3[9760]<=16'd23752; ROM4[9760]<=16'd57228;
ROM1[9761]<=16'd4795; ROM2[9761]<=16'd0; ROM3[9761]<=16'd23771; ROM4[9761]<=16'd57245;
ROM1[9762]<=16'd4794; ROM2[9762]<=16'd0; ROM3[9762]<=16'd23763; ROM4[9762]<=16'd57243;
ROM1[9763]<=16'd4791; ROM2[9763]<=16'd0; ROM3[9763]<=16'd23725; ROM4[9763]<=16'd57213;
ROM1[9764]<=16'd4828; ROM2[9764]<=16'd0; ROM3[9764]<=16'd23716; ROM4[9764]<=16'd57214;
ROM1[9765]<=16'd4845; ROM2[9765]<=16'd0; ROM3[9765]<=16'd23714; ROM4[9765]<=16'd57218;
ROM1[9766]<=16'd4836; ROM2[9766]<=16'd0; ROM3[9766]<=16'd23719; ROM4[9766]<=16'd57218;
ROM1[9767]<=16'd4836; ROM2[9767]<=16'd0; ROM3[9767]<=16'd23741; ROM4[9767]<=16'd57234;
ROM1[9768]<=16'd4830; ROM2[9768]<=16'd0; ROM3[9768]<=16'd23748; ROM4[9768]<=16'd57239;
ROM1[9769]<=16'd4802; ROM2[9769]<=16'd0; ROM3[9769]<=16'd23739; ROM4[9769]<=16'd57225;
ROM1[9770]<=16'd4794; ROM2[9770]<=16'd0; ROM3[9770]<=16'd23738; ROM4[9770]<=16'd57220;
ROM1[9771]<=16'd4816; ROM2[9771]<=16'd0; ROM3[9771]<=16'd23738; ROM4[9771]<=16'd57224;
ROM1[9772]<=16'd4846; ROM2[9772]<=16'd0; ROM3[9772]<=16'd23723; ROM4[9772]<=16'd57220;
ROM1[9773]<=16'd4870; ROM2[9773]<=16'd0; ROM3[9773]<=16'd23715; ROM4[9773]<=16'd57222;
ROM1[9774]<=16'd4879; ROM2[9774]<=16'd0; ROM3[9774]<=16'd23737; ROM4[9774]<=16'd57243;
ROM1[9775]<=16'd4889; ROM2[9775]<=16'd0; ROM3[9775]<=16'd23773; ROM4[9775]<=16'd57275;
ROM1[9776]<=16'd4854; ROM2[9776]<=16'd0; ROM3[9776]<=16'd23760; ROM4[9776]<=16'd57254;
ROM1[9777]<=16'd4813; ROM2[9777]<=16'd0; ROM3[9777]<=16'd23741; ROM4[9777]<=16'd57225;
ROM1[9778]<=16'd4811; ROM2[9778]<=16'd0; ROM3[9778]<=16'd23744; ROM4[9778]<=16'd57229;
ROM1[9779]<=16'd4790; ROM2[9779]<=16'd0; ROM3[9779]<=16'd23716; ROM4[9779]<=16'd57204;
ROM1[9780]<=16'd4822; ROM2[9780]<=16'd0; ROM3[9780]<=16'd23720; ROM4[9780]<=16'd57215;
ROM1[9781]<=16'd4864; ROM2[9781]<=16'd0; ROM3[9781]<=16'd23725; ROM4[9781]<=16'd57231;
ROM1[9782]<=16'd4837; ROM2[9782]<=16'd0; ROM3[9782]<=16'd23700; ROM4[9782]<=16'd57203;
ROM1[9783]<=16'd4805; ROM2[9783]<=16'd0; ROM3[9783]<=16'd23690; ROM4[9783]<=16'd57186;
ROM1[9784]<=16'd4784; ROM2[9784]<=16'd0; ROM3[9784]<=16'd23695; ROM4[9784]<=16'd57183;
ROM1[9785]<=16'd4777; ROM2[9785]<=16'd0; ROM3[9785]<=16'd23705; ROM4[9785]<=16'd57191;
ROM1[9786]<=16'd4766; ROM2[9786]<=16'd0; ROM3[9786]<=16'd23712; ROM4[9786]<=16'd57197;
ROM1[9787]<=16'd4778; ROM2[9787]<=16'd0; ROM3[9787]<=16'd23726; ROM4[9787]<=16'd57208;
ROM1[9788]<=16'd4793; ROM2[9788]<=16'd0; ROM3[9788]<=16'd23715; ROM4[9788]<=16'd57203;
ROM1[9789]<=16'd4813; ROM2[9789]<=16'd0; ROM3[9789]<=16'd23696; ROM4[9789]<=16'd57196;
ROM1[9790]<=16'd4824; ROM2[9790]<=16'd0; ROM3[9790]<=16'd23695; ROM4[9790]<=16'd57198;
ROM1[9791]<=16'd4807; ROM2[9791]<=16'd0; ROM3[9791]<=16'd23702; ROM4[9791]<=16'd57198;
ROM1[9792]<=16'd4788; ROM2[9792]<=16'd0; ROM3[9792]<=16'd23716; ROM4[9792]<=16'd57204;
ROM1[9793]<=16'd4773; ROM2[9793]<=16'd0; ROM3[9793]<=16'd23721; ROM4[9793]<=16'd57205;
ROM1[9794]<=16'd4751; ROM2[9794]<=16'd0; ROM3[9794]<=16'd23722; ROM4[9794]<=16'd57201;
ROM1[9795]<=16'd4740; ROM2[9795]<=16'd0; ROM3[9795]<=16'd23725; ROM4[9795]<=16'd57200;
ROM1[9796]<=16'd4752; ROM2[9796]<=16'd0; ROM3[9796]<=16'd23720; ROM4[9796]<=16'd57204;
ROM1[9797]<=16'd4786; ROM2[9797]<=16'd0; ROM3[9797]<=16'd23712; ROM4[9797]<=16'd57207;
ROM1[9798]<=16'd4807; ROM2[9798]<=16'd0; ROM3[9798]<=16'd23701; ROM4[9798]<=16'd57205;
ROM1[9799]<=16'd4799; ROM2[9799]<=16'd0; ROM3[9799]<=16'd23700; ROM4[9799]<=16'd57205;
ROM1[9800]<=16'd4784; ROM2[9800]<=16'd0; ROM3[9800]<=16'd23711; ROM4[9800]<=16'd57207;
ROM1[9801]<=16'd4772; ROM2[9801]<=16'd0; ROM3[9801]<=16'd23729; ROM4[9801]<=16'd57214;
ROM1[9802]<=16'd4760; ROM2[9802]<=16'd0; ROM3[9802]<=16'd23742; ROM4[9802]<=16'd57220;
ROM1[9803]<=16'd4759; ROM2[9803]<=16'd0; ROM3[9803]<=16'd23749; ROM4[9803]<=16'd57228;
ROM1[9804]<=16'd4773; ROM2[9804]<=16'd0; ROM3[9804]<=16'd23753; ROM4[9804]<=16'd57234;
ROM1[9805]<=16'd4799; ROM2[9805]<=16'd0; ROM3[9805]<=16'd23749; ROM4[9805]<=16'd57239;
ROM1[9806]<=16'd4825; ROM2[9806]<=16'd0; ROM3[9806]<=16'd23734; ROM4[9806]<=16'd57235;
ROM1[9807]<=16'd4825; ROM2[9807]<=16'd0; ROM3[9807]<=16'd23733; ROM4[9807]<=16'd57235;
ROM1[9808]<=16'd4825; ROM2[9808]<=16'd0; ROM3[9808]<=16'd23759; ROM4[9808]<=16'd57253;
ROM1[9809]<=16'd4815; ROM2[9809]<=16'd0; ROM3[9809]<=16'd23775; ROM4[9809]<=16'd57257;
ROM1[9810]<=16'd4792; ROM2[9810]<=16'd0; ROM3[9810]<=16'd23768; ROM4[9810]<=16'd57245;
ROM1[9811]<=16'd4787; ROM2[9811]<=16'd0; ROM3[9811]<=16'd23775; ROM4[9811]<=16'd57249;
ROM1[9812]<=16'd4785; ROM2[9812]<=16'd0; ROM3[9812]<=16'd23766; ROM4[9812]<=16'd57243;
ROM1[9813]<=16'd4773; ROM2[9813]<=16'd0; ROM3[9813]<=16'd23723; ROM4[9813]<=16'd57211;
ROM1[9814]<=16'd4802; ROM2[9814]<=16'd0; ROM3[9814]<=16'd23706; ROM4[9814]<=16'd57205;
ROM1[9815]<=16'd4817; ROM2[9815]<=16'd0; ROM3[9815]<=16'd23706; ROM4[9815]<=16'd57208;
ROM1[9816]<=16'd4809; ROM2[9816]<=16'd0; ROM3[9816]<=16'd23713; ROM4[9816]<=16'd57214;
ROM1[9817]<=16'd4806; ROM2[9817]<=16'd0; ROM3[9817]<=16'd23730; ROM4[9817]<=16'd57226;
ROM1[9818]<=16'd4790; ROM2[9818]<=16'd0; ROM3[9818]<=16'd23732; ROM4[9818]<=16'd57219;
ROM1[9819]<=16'd4752; ROM2[9819]<=16'd0; ROM3[9819]<=16'd23707; ROM4[9819]<=16'd57189;
ROM1[9820]<=16'd4740; ROM2[9820]<=16'd0; ROM3[9820]<=16'd23691; ROM4[9820]<=16'd57168;
ROM1[9821]<=16'd4763; ROM2[9821]<=16'd0; ROM3[9821]<=16'd23693; ROM4[9821]<=16'd57175;
ROM1[9822]<=16'd4796; ROM2[9822]<=16'd0; ROM3[9822]<=16'd23688; ROM4[9822]<=16'd57181;
ROM1[9823]<=16'd4818; ROM2[9823]<=16'd0; ROM3[9823]<=16'd23687; ROM4[9823]<=16'd57184;
ROM1[9824]<=16'd4804; ROM2[9824]<=16'd0; ROM3[9824]<=16'd23686; ROM4[9824]<=16'd57178;
ROM1[9825]<=16'd4781; ROM2[9825]<=16'd0; ROM3[9825]<=16'd23691; ROM4[9825]<=16'd57175;
ROM1[9826]<=16'd4775; ROM2[9826]<=16'd0; ROM3[9826]<=16'd23706; ROM4[9826]<=16'd57184;
ROM1[9827]<=16'd4767; ROM2[9827]<=16'd0; ROM3[9827]<=16'd23715; ROM4[9827]<=16'd57191;
ROM1[9828]<=16'd4759; ROM2[9828]<=16'd0; ROM3[9828]<=16'd23723; ROM4[9828]<=16'd57194;
ROM1[9829]<=16'd4784; ROM2[9829]<=16'd0; ROM3[9829]<=16'd23735; ROM4[9829]<=16'd57207;
ROM1[9830]<=16'd4824; ROM2[9830]<=16'd0; ROM3[9830]<=16'd23738; ROM4[9830]<=16'd57217;
ROM1[9831]<=16'd4853; ROM2[9831]<=16'd0; ROM3[9831]<=16'd23731; ROM4[9831]<=16'd57219;
ROM1[9832]<=16'd4850; ROM2[9832]<=16'd0; ROM3[9832]<=16'd23730; ROM4[9832]<=16'd57219;
ROM1[9833]<=16'd4816; ROM2[9833]<=16'd0; ROM3[9833]<=16'd23724; ROM4[9833]<=16'd57203;
ROM1[9834]<=16'd4788; ROM2[9834]<=16'd0; ROM3[9834]<=16'd23726; ROM4[9834]<=16'd57194;
ROM1[9835]<=16'd4783; ROM2[9835]<=16'd0; ROM3[9835]<=16'd23739; ROM4[9835]<=16'd57202;
ROM1[9836]<=16'd4768; ROM2[9836]<=16'd0; ROM3[9836]<=16'd23747; ROM4[9836]<=16'd57207;
ROM1[9837]<=16'd4768; ROM2[9837]<=16'd0; ROM3[9837]<=16'd23749; ROM4[9837]<=16'd57212;
ROM1[9838]<=16'd4785; ROM2[9838]<=16'd0; ROM3[9838]<=16'd23739; ROM4[9838]<=16'd57212;
ROM1[9839]<=16'd4803; ROM2[9839]<=16'd0; ROM3[9839]<=16'd23716; ROM4[9839]<=16'd57199;
ROM1[9840]<=16'd4807; ROM2[9840]<=16'd0; ROM3[9840]<=16'd23707; ROM4[9840]<=16'd57191;
ROM1[9841]<=16'd4791; ROM2[9841]<=16'd0; ROM3[9841]<=16'd23717; ROM4[9841]<=16'd57195;
ROM1[9842]<=16'd4777; ROM2[9842]<=16'd0; ROM3[9842]<=16'd23737; ROM4[9842]<=16'd57201;
ROM1[9843]<=16'd4776; ROM2[9843]<=16'd0; ROM3[9843]<=16'd23751; ROM4[9843]<=16'd57205;
ROM1[9844]<=16'd4761; ROM2[9844]<=16'd0; ROM3[9844]<=16'd23755; ROM4[9844]<=16'd57208;
ROM1[9845]<=16'd4756; ROM2[9845]<=16'd0; ROM3[9845]<=16'd23756; ROM4[9845]<=16'd57206;
ROM1[9846]<=16'd4784; ROM2[9846]<=16'd0; ROM3[9846]<=16'd23762; ROM4[9846]<=16'd57219;
ROM1[9847]<=16'd4800; ROM2[9847]<=16'd0; ROM3[9847]<=16'd23745; ROM4[9847]<=16'd57217;
ROM1[9848]<=16'd4800; ROM2[9848]<=16'd0; ROM3[9848]<=16'd23722; ROM4[9848]<=16'd57195;
ROM1[9849]<=16'd4796; ROM2[9849]<=16'd0; ROM3[9849]<=16'd23727; ROM4[9849]<=16'd57194;
ROM1[9850]<=16'd4780; ROM2[9850]<=16'd0; ROM3[9850]<=16'd23733; ROM4[9850]<=16'd57195;
ROM1[9851]<=16'd4769; ROM2[9851]<=16'd0; ROM3[9851]<=16'd23746; ROM4[9851]<=16'd57200;
ROM1[9852]<=16'd4766; ROM2[9852]<=16'd0; ROM3[9852]<=16'd23761; ROM4[9852]<=16'd57212;
ROM1[9853]<=16'd4749; ROM2[9853]<=16'd0; ROM3[9853]<=16'd23758; ROM4[9853]<=16'd57203;
ROM1[9854]<=16'd4742; ROM2[9854]<=16'd0; ROM3[9854]<=16'd23747; ROM4[9854]<=16'd57194;
ROM1[9855]<=16'd4769; ROM2[9855]<=16'd0; ROM3[9855]<=16'd23740; ROM4[9855]<=16'd57194;
ROM1[9856]<=16'd4810; ROM2[9856]<=16'd0; ROM3[9856]<=16'd23739; ROM4[9856]<=16'd57203;
ROM1[9857]<=16'd4825; ROM2[9857]<=16'd0; ROM3[9857]<=16'd23748; ROM4[9857]<=16'd57218;
ROM1[9858]<=16'd4802; ROM2[9858]<=16'd0; ROM3[9858]<=16'd23743; ROM4[9858]<=16'd57208;
ROM1[9859]<=16'd4773; ROM2[9859]<=16'd0; ROM3[9859]<=16'd23738; ROM4[9859]<=16'd57199;
ROM1[9860]<=16'd4754; ROM2[9860]<=16'd0; ROM3[9860]<=16'd23733; ROM4[9860]<=16'd57193;
ROM1[9861]<=16'd4725; ROM2[9861]<=16'd0; ROM3[9861]<=16'd23725; ROM4[9861]<=16'd57179;
ROM1[9862]<=16'd4729; ROM2[9862]<=16'd0; ROM3[9862]<=16'd23730; ROM4[9862]<=16'd57180;
ROM1[9863]<=16'd4764; ROM2[9863]<=16'd0; ROM3[9863]<=16'd23731; ROM4[9863]<=16'd57189;
ROM1[9864]<=16'd4813; ROM2[9864]<=16'd0; ROM3[9864]<=16'd23735; ROM4[9864]<=16'd57206;
ROM1[9865]<=16'd4840; ROM2[9865]<=16'd0; ROM3[9865]<=16'd23745; ROM4[9865]<=16'd57221;
ROM1[9866]<=16'd4818; ROM2[9866]<=16'd0; ROM3[9866]<=16'd23746; ROM4[9866]<=16'd57216;
ROM1[9867]<=16'd4788; ROM2[9867]<=16'd0; ROM3[9867]<=16'd23746; ROM4[9867]<=16'd57209;
ROM1[9868]<=16'd4770; ROM2[9868]<=16'd0; ROM3[9868]<=16'd23749; ROM4[9868]<=16'd57202;
ROM1[9869]<=16'd4760; ROM2[9869]<=16'd0; ROM3[9869]<=16'd23760; ROM4[9869]<=16'd57206;
ROM1[9870]<=16'd4757; ROM2[9870]<=16'd0; ROM3[9870]<=16'd23760; ROM4[9870]<=16'd57208;
ROM1[9871]<=16'd4764; ROM2[9871]<=16'd0; ROM3[9871]<=16'd23746; ROM4[9871]<=16'd57199;
ROM1[9872]<=16'd4788; ROM2[9872]<=16'd0; ROM3[9872]<=16'd23729; ROM4[9872]<=16'd57194;
ROM1[9873]<=16'd4799; ROM2[9873]<=16'd0; ROM3[9873]<=16'd23711; ROM4[9873]<=16'd57190;
ROM1[9874]<=16'd4795; ROM2[9874]<=16'd0; ROM3[9874]<=16'd23721; ROM4[9874]<=16'd57201;
ROM1[9875]<=16'd4787; ROM2[9875]<=16'd0; ROM3[9875]<=16'd23741; ROM4[9875]<=16'd57212;
ROM1[9876]<=16'd4771; ROM2[9876]<=16'd0; ROM3[9876]<=16'd23750; ROM4[9876]<=16'd57211;
ROM1[9877]<=16'd4745; ROM2[9877]<=16'd0; ROM3[9877]<=16'd23749; ROM4[9877]<=16'd57203;
ROM1[9878]<=16'd4734; ROM2[9878]<=16'd0; ROM3[9878]<=16'd23750; ROM4[9878]<=16'd57202;
ROM1[9879]<=16'd4743; ROM2[9879]<=16'd0; ROM3[9879]<=16'd23752; ROM4[9879]<=16'd57205;
ROM1[9880]<=16'd4766; ROM2[9880]<=16'd0; ROM3[9880]<=16'd23740; ROM4[9880]<=16'd57202;
ROM1[9881]<=16'd4799; ROM2[9881]<=16'd0; ROM3[9881]<=16'd23728; ROM4[9881]<=16'd57203;
ROM1[9882]<=16'd4807; ROM2[9882]<=16'd0; ROM3[9882]<=16'd23738; ROM4[9882]<=16'd57215;
ROM1[9883]<=16'd4794; ROM2[9883]<=16'd0; ROM3[9883]<=16'd23752; ROM4[9883]<=16'd57222;
ROM1[9884]<=16'd4790; ROM2[9884]<=16'd0; ROM3[9884]<=16'd23775; ROM4[9884]<=16'd57239;
ROM1[9885]<=16'd4785; ROM2[9885]<=16'd0; ROM3[9885]<=16'd23787; ROM4[9885]<=16'd57246;
ROM1[9886]<=16'd4756; ROM2[9886]<=16'd0; ROM3[9886]<=16'd23772; ROM4[9886]<=16'd57225;
ROM1[9887]<=16'd4750; ROM2[9887]<=16'd0; ROM3[9887]<=16'd23764; ROM4[9887]<=16'd57218;
ROM1[9888]<=16'd4765; ROM2[9888]<=16'd0; ROM3[9888]<=16'd23754; ROM4[9888]<=16'd57217;
ROM1[9889]<=16'd4798; ROM2[9889]<=16'd0; ROM3[9889]<=16'd23742; ROM4[9889]<=16'd57214;
ROM1[9890]<=16'd4820; ROM2[9890]<=16'd0; ROM3[9890]<=16'd23743; ROM4[9890]<=16'd57223;
ROM1[9891]<=16'd4809; ROM2[9891]<=16'd0; ROM3[9891]<=16'd23751; ROM4[9891]<=16'd57231;
ROM1[9892]<=16'd4792; ROM2[9892]<=16'd0; ROM3[9892]<=16'd23761; ROM4[9892]<=16'd57231;
ROM1[9893]<=16'd4781; ROM2[9893]<=16'd0; ROM3[9893]<=16'd23767; ROM4[9893]<=16'd57231;
ROM1[9894]<=16'd4770; ROM2[9894]<=16'd0; ROM3[9894]<=16'd23772; ROM4[9894]<=16'd57231;
ROM1[9895]<=16'd4770; ROM2[9895]<=16'd0; ROM3[9895]<=16'd23777; ROM4[9895]<=16'd57233;
ROM1[9896]<=16'd4786; ROM2[9896]<=16'd0; ROM3[9896]<=16'd23765; ROM4[9896]<=16'd57228;
ROM1[9897]<=16'd4802; ROM2[9897]<=16'd0; ROM3[9897]<=16'd23745; ROM4[9897]<=16'd57218;
ROM1[9898]<=16'd4815; ROM2[9898]<=16'd0; ROM3[9898]<=16'd23728; ROM4[9898]<=16'd57207;
ROM1[9899]<=16'd4803; ROM2[9899]<=16'd0; ROM3[9899]<=16'd23723; ROM4[9899]<=16'd57199;
ROM1[9900]<=16'd4787; ROM2[9900]<=16'd0; ROM3[9900]<=16'd23733; ROM4[9900]<=16'd57202;
ROM1[9901]<=16'd4776; ROM2[9901]<=16'd0; ROM3[9901]<=16'd23739; ROM4[9901]<=16'd57202;
ROM1[9902]<=16'd4768; ROM2[9902]<=16'd0; ROM3[9902]<=16'd23750; ROM4[9902]<=16'd57207;
ROM1[9903]<=16'd4764; ROM2[9903]<=16'd0; ROM3[9903]<=16'd23760; ROM4[9903]<=16'd57214;
ROM1[9904]<=16'd4769; ROM2[9904]<=16'd0; ROM3[9904]<=16'd23759; ROM4[9904]<=16'd57213;
ROM1[9905]<=16'd4781; ROM2[9905]<=16'd0; ROM3[9905]<=16'd23742; ROM4[9905]<=16'd57205;
ROM1[9906]<=16'd4808; ROM2[9906]<=16'd0; ROM3[9906]<=16'd23729; ROM4[9906]<=16'd57202;
ROM1[9907]<=16'd4814; ROM2[9907]<=16'd0; ROM3[9907]<=16'd23734; ROM4[9907]<=16'd57207;
ROM1[9908]<=16'd4801; ROM2[9908]<=16'd0; ROM3[9908]<=16'd23737; ROM4[9908]<=16'd57204;
ROM1[9909]<=16'd4819; ROM2[9909]<=16'd0; ROM3[9909]<=16'd23771; ROM4[9909]<=16'd57236;
ROM1[9910]<=16'd4823; ROM2[9910]<=16'd0; ROM3[9910]<=16'd23791; ROM4[9910]<=16'd57249;
ROM1[9911]<=16'd4796; ROM2[9911]<=16'd0; ROM3[9911]<=16'd23780; ROM4[9911]<=16'd57232;
ROM1[9912]<=16'd4774; ROM2[9912]<=16'd0; ROM3[9912]<=16'd23755; ROM4[9912]<=16'd57210;
ROM1[9913]<=16'd4771; ROM2[9913]<=16'd0; ROM3[9913]<=16'd23727; ROM4[9913]<=16'd57186;
ROM1[9914]<=16'd4797; ROM2[9914]<=16'd0; ROM3[9914]<=16'd23713; ROM4[9914]<=16'd57184;
ROM1[9915]<=16'd4818; ROM2[9915]<=16'd0; ROM3[9915]<=16'd23715; ROM4[9915]<=16'd57191;
ROM1[9916]<=16'd4828; ROM2[9916]<=16'd0; ROM3[9916]<=16'd23745; ROM4[9916]<=16'd57210;
ROM1[9917]<=16'd4807; ROM2[9917]<=16'd0; ROM3[9917]<=16'd23752; ROM4[9917]<=16'd57211;
ROM1[9918]<=16'd4784; ROM2[9918]<=16'd0; ROM3[9918]<=16'd23745; ROM4[9918]<=16'd57203;
ROM1[9919]<=16'd4767; ROM2[9919]<=16'd0; ROM3[9919]<=16'd23750; ROM4[9919]<=16'd57202;
ROM1[9920]<=16'd4748; ROM2[9920]<=16'd0; ROM3[9920]<=16'd23742; ROM4[9920]<=16'd57192;
ROM1[9921]<=16'd4757; ROM2[9921]<=16'd0; ROM3[9921]<=16'd23734; ROM4[9921]<=16'd57186;
ROM1[9922]<=16'd4790; ROM2[9922]<=16'd0; ROM3[9922]<=16'd23728; ROM4[9922]<=16'd57188;
ROM1[9923]<=16'd4810; ROM2[9923]<=16'd0; ROM3[9923]<=16'd23719; ROM4[9923]<=16'd57191;
ROM1[9924]<=16'd4821; ROM2[9924]<=16'd0; ROM3[9924]<=16'd23735; ROM4[9924]<=16'd57209;
ROM1[9925]<=16'd4809; ROM2[9925]<=16'd0; ROM3[9925]<=16'd23744; ROM4[9925]<=16'd57213;
ROM1[9926]<=16'd4771; ROM2[9926]<=16'd0; ROM3[9926]<=16'd23734; ROM4[9926]<=16'd57190;
ROM1[9927]<=16'd4757; ROM2[9927]<=16'd0; ROM3[9927]<=16'd23739; ROM4[9927]<=16'd57188;
ROM1[9928]<=16'd4750; ROM2[9928]<=16'd0; ROM3[9928]<=16'd23740; ROM4[9928]<=16'd57189;
ROM1[9929]<=16'd4758; ROM2[9929]<=16'd0; ROM3[9929]<=16'd23745; ROM4[9929]<=16'd57193;
ROM1[9930]<=16'd4804; ROM2[9930]<=16'd0; ROM3[9930]<=16'd23756; ROM4[9930]<=16'd57215;
ROM1[9931]<=16'd4836; ROM2[9931]<=16'd0; ROM3[9931]<=16'd23747; ROM4[9931]<=16'd57219;
ROM1[9932]<=16'd4826; ROM2[9932]<=16'd0; ROM3[9932]<=16'd23739; ROM4[9932]<=16'd57210;
ROM1[9933]<=16'd4803; ROM2[9933]<=16'd0; ROM3[9933]<=16'd23739; ROM4[9933]<=16'd57205;
ROM1[9934]<=16'd4781; ROM2[9934]<=16'd0; ROM3[9934]<=16'd23741; ROM4[9934]<=16'd57202;
ROM1[9935]<=16'd4769; ROM2[9935]<=16'd0; ROM3[9935]<=16'd23752; ROM4[9935]<=16'd57202;
ROM1[9936]<=16'd4761; ROM2[9936]<=16'd0; ROM3[9936]<=16'd23760; ROM4[9936]<=16'd57205;
ROM1[9937]<=16'd4770; ROM2[9937]<=16'd0; ROM3[9937]<=16'd23765; ROM4[9937]<=16'd57210;
ROM1[9938]<=16'd4795; ROM2[9938]<=16'd0; ROM3[9938]<=16'd23760; ROM4[9938]<=16'd57215;
ROM1[9939]<=16'd4822; ROM2[9939]<=16'd0; ROM3[9939]<=16'd23746; ROM4[9939]<=16'd57212;
ROM1[9940]<=16'd4828; ROM2[9940]<=16'd0; ROM3[9940]<=16'd23740; ROM4[9940]<=16'd57206;
ROM1[9941]<=16'd4825; ROM2[9941]<=16'd0; ROM3[9941]<=16'd23757; ROM4[9941]<=16'd57217;
ROM1[9942]<=16'd4829; ROM2[9942]<=16'd0; ROM3[9942]<=16'd23782; ROM4[9942]<=16'd57237;
ROM1[9943]<=16'd4806; ROM2[9943]<=16'd0; ROM3[9943]<=16'd23771; ROM4[9943]<=16'd57226;
ROM1[9944]<=16'd4775; ROM2[9944]<=16'd0; ROM3[9944]<=16'd23757; ROM4[9944]<=16'd57214;
ROM1[9945]<=16'd4775; ROM2[9945]<=16'd0; ROM3[9945]<=16'd23759; ROM4[9945]<=16'd57217;
ROM1[9946]<=16'd4780; ROM2[9946]<=16'd0; ROM3[9946]<=16'd23747; ROM4[9946]<=16'd57208;
ROM1[9947]<=16'd4819; ROM2[9947]<=16'd0; ROM3[9947]<=16'd23746; ROM4[9947]<=16'd57218;
ROM1[9948]<=16'd4849; ROM2[9948]<=16'd0; ROM3[9948]<=16'd23742; ROM4[9948]<=16'd57221;
ROM1[9949]<=16'd4835; ROM2[9949]<=16'd0; ROM3[9949]<=16'd23730; ROM4[9949]<=16'd57212;
ROM1[9950]<=16'd4814; ROM2[9950]<=16'd0; ROM3[9950]<=16'd23736; ROM4[9950]<=16'd57215;
ROM1[9951]<=16'd4809; ROM2[9951]<=16'd0; ROM3[9951]<=16'd23755; ROM4[9951]<=16'd57224;
ROM1[9952]<=16'd4799; ROM2[9952]<=16'd0; ROM3[9952]<=16'd23762; ROM4[9952]<=16'd57222;
ROM1[9953]<=16'd4774; ROM2[9953]<=16'd0; ROM3[9953]<=16'd23758; ROM4[9953]<=16'd57215;
ROM1[9954]<=16'd4776; ROM2[9954]<=16'd0; ROM3[9954]<=16'd23759; ROM4[9954]<=16'd57212;
ROM1[9955]<=16'd4812; ROM2[9955]<=16'd0; ROM3[9955]<=16'd23761; ROM4[9955]<=16'd57222;
ROM1[9956]<=16'd4859; ROM2[9956]<=16'd0; ROM3[9956]<=16'd23774; ROM4[9956]<=16'd57248;
ROM1[9957]<=16'd4880; ROM2[9957]<=16'd0; ROM3[9957]<=16'd23799; ROM4[9957]<=16'd57271;
ROM1[9958]<=16'd4854; ROM2[9958]<=16'd0; ROM3[9958]<=16'd23792; ROM4[9958]<=16'd57260;
ROM1[9959]<=16'd4805; ROM2[9959]<=16'd0; ROM3[9959]<=16'd23771; ROM4[9959]<=16'd57234;
ROM1[9960]<=16'd4789; ROM2[9960]<=16'd0; ROM3[9960]<=16'd23779; ROM4[9960]<=16'd57239;
ROM1[9961]<=16'd4775; ROM2[9961]<=16'd0; ROM3[9961]<=16'd23785; ROM4[9961]<=16'd57236;
ROM1[9962]<=16'd4786; ROM2[9962]<=16'd0; ROM3[9962]<=16'd23796; ROM4[9962]<=16'd57242;
ROM1[9963]<=16'd4818; ROM2[9963]<=16'd0; ROM3[9963]<=16'd23799; ROM4[9963]<=16'd57252;
ROM1[9964]<=16'd4821; ROM2[9964]<=16'd0; ROM3[9964]<=16'd23755; ROM4[9964]<=16'd57223;
ROM1[9965]<=16'd4812; ROM2[9965]<=16'd0; ROM3[9965]<=16'd23731; ROM4[9965]<=16'd57206;
ROM1[9966]<=16'd4803; ROM2[9966]<=16'd0; ROM3[9966]<=16'd23744; ROM4[9966]<=16'd57210;
ROM1[9967]<=16'd4794; ROM2[9967]<=16'd0; ROM3[9967]<=16'd23757; ROM4[9967]<=16'd57218;
ROM1[9968]<=16'd4799; ROM2[9968]<=16'd0; ROM3[9968]<=16'd23778; ROM4[9968]<=16'd57229;
ROM1[9969]<=16'd4792; ROM2[9969]<=16'd0; ROM3[9969]<=16'd23785; ROM4[9969]<=16'd57230;
ROM1[9970]<=16'd4776; ROM2[9970]<=16'd0; ROM3[9970]<=16'd23772; ROM4[9970]<=16'd57221;
ROM1[9971]<=16'd4791; ROM2[9971]<=16'd0; ROM3[9971]<=16'd23762; ROM4[9971]<=16'd57220;
ROM1[9972]<=16'd4819; ROM2[9972]<=16'd0; ROM3[9972]<=16'd23746; ROM4[9972]<=16'd57218;
ROM1[9973]<=16'd4842; ROM2[9973]<=16'd0; ROM3[9973]<=16'd23745; ROM4[9973]<=16'd57225;
ROM1[9974]<=16'd4844; ROM2[9974]<=16'd0; ROM3[9974]<=16'd23754; ROM4[9974]<=16'd57235;
ROM1[9975]<=16'd4819; ROM2[9975]<=16'd0; ROM3[9975]<=16'd23761; ROM4[9975]<=16'd57229;
ROM1[9976]<=16'd4799; ROM2[9976]<=16'd0; ROM3[9976]<=16'd23771; ROM4[9976]<=16'd57228;
ROM1[9977]<=16'd4776; ROM2[9977]<=16'd0; ROM3[9977]<=16'd23764; ROM4[9977]<=16'd57221;
ROM1[9978]<=16'd4761; ROM2[9978]<=16'd0; ROM3[9978]<=16'd23759; ROM4[9978]<=16'd57214;
ROM1[9979]<=16'd4778; ROM2[9979]<=16'd0; ROM3[9979]<=16'd23764; ROM4[9979]<=16'd57223;
ROM1[9980]<=16'd4805; ROM2[9980]<=16'd0; ROM3[9980]<=16'd23755; ROM4[9980]<=16'd57223;
ROM1[9981]<=16'd4815; ROM2[9981]<=16'd0; ROM3[9981]<=16'd23722; ROM4[9981]<=16'd57203;
ROM1[9982]<=16'd4809; ROM2[9982]<=16'd0; ROM3[9982]<=16'd23716; ROM4[9982]<=16'd57198;
ROM1[9983]<=16'd4790; ROM2[9983]<=16'd0; ROM3[9983]<=16'd23715; ROM4[9983]<=16'd57190;
ROM1[9984]<=16'd4772; ROM2[9984]<=16'd0; ROM3[9984]<=16'd23718; ROM4[9984]<=16'd57184;
ROM1[9985]<=16'd4774; ROM2[9985]<=16'd0; ROM3[9985]<=16'd23732; ROM4[9985]<=16'd57195;
ROM1[9986]<=16'd4774; ROM2[9986]<=16'd0; ROM3[9986]<=16'd23746; ROM4[9986]<=16'd57206;
ROM1[9987]<=16'd4785; ROM2[9987]<=16'd0; ROM3[9987]<=16'd23752; ROM4[9987]<=16'd57214;
ROM1[9988]<=16'd4792; ROM2[9988]<=16'd0; ROM3[9988]<=16'd23730; ROM4[9988]<=16'd57199;
ROM1[9989]<=16'd4828; ROM2[9989]<=16'd0; ROM3[9989]<=16'd23722; ROM4[9989]<=16'd57204;
ROM1[9990]<=16'd4844; ROM2[9990]<=16'd0; ROM3[9990]<=16'd23719; ROM4[9990]<=16'd57206;
ROM1[9991]<=16'd4816; ROM2[9991]<=16'd0; ROM3[9991]<=16'd23709; ROM4[9991]<=16'd57197;
ROM1[9992]<=16'd4804; ROM2[9992]<=16'd0; ROM3[9992]<=16'd23725; ROM4[9992]<=16'd57206;
ROM1[9993]<=16'd4801; ROM2[9993]<=16'd0; ROM3[9993]<=16'd23744; ROM4[9993]<=16'd57215;
ROM1[9994]<=16'd4783; ROM2[9994]<=16'd0; ROM3[9994]<=16'd23748; ROM4[9994]<=16'd57213;
ROM1[9995]<=16'd4776; ROM2[9995]<=16'd0; ROM3[9995]<=16'd23746; ROM4[9995]<=16'd57207;
ROM1[9996]<=16'd4795; ROM2[9996]<=16'd0; ROM3[9996]<=16'd23747; ROM4[9996]<=16'd57215;
ROM1[9997]<=16'd4828; ROM2[9997]<=16'd0; ROM3[9997]<=16'd23744; ROM4[9997]<=16'd57223;
ROM1[9998]<=16'd4854; ROM2[9998]<=16'd0; ROM3[9998]<=16'd23740; ROM4[9998]<=16'd57228;
ROM1[9999]<=16'd4848; ROM2[9999]<=16'd0; ROM3[9999]<=16'd23747; ROM4[9999]<=16'd57229;
	end
	else begin
		if(cnt == 127) begin
				cnt<=0;
			end
		//원래는 addr이다.
		data1 <= ROM1[cnt];
		data2 <= ROM2[cnt];
		data3 <= ROM3[cnt];
		data4 <= ROM4[cnt];
		cnt <= cnt+1;
	end
end
endmodule 
